`timescale 1ns / 1ps
`include "defines.vh"

module encoder
(
    input wire [31:0] data,
    output reg [4:0] code
);

always @(*)
begin
    casez (data)
        // 从最高位(31)到最低位(0)的优先级顺序
        32'b1???????_????????_????????_????????: code = 5'd31;  // 位31
        32'b01??????_????????_????????_????????: code = 5'd30;  // 位30
        32'b001?????_????????_????????_????????: code = 5'd29;  // 位29
        32'b0001????_????????_????????_????????: code = 5'd28;  // 位28
        32'b00001???_????????_????????_????????: code = 5'd27;  // 位27
        32'b000001??_????????_????????_????????: code = 5'd26;  // 位26
        32'b0000001?_????????_????????_????????: code = 5'd25;  // 位25
        32'b00000001_????????_????????_????????: code = 5'd24;  // 位24
        32'b00000000_1???????_????????_????????: code = 5'd23;  // 位23
        32'b00000000_01??????_????????_????????: code = 5'd22;  // 位22
        32'b00000000_001?????_????????_????????: code = 5'd21;  // 位21
        32'b00000000_0001????_????????_????????: code = 5'd20;  // 位20
        32'b00000000_00001???_????????_????????: code = 5'd19;  // 位19
        32'b00000000_000001??_????????_????????: code = 5'd18;  // 位18
        32'b00000000_0000001?_????????_????????: code = 5'd17;  // 位17
        32'b00000000_00000001_????????_????????: code = 5'd16;  // 位16
        32'b00000000_00000000_1???????_????????: code = 5'd15;  // 位15
        32'b00000000_00000000_01??????_????????: code = 5'd14;  // 位14
        32'b00000000_00000000_001?????_????????: code = 5'd13;  // 位13
        32'b00000000_00000000_0001????_????????: code = 5'd12;  // 位12
        32'b00000000_00000000_00001???_????????: code = 5'd11;  // 位11
        32'b00000000_00000000_000001??_????????: code = 5'd10;  // 位10
        32'b00000000_00000000_0000001?_????????: code = 5'd9;   // 位9
        32'b00000000_00000000_00000001_????????: code = 5'd8;   // 位8
        32'b00000000_00000000_00000000_1???????: code = 5'd7;   // 位7
        32'b00000000_00000000_00000000_01??????: code = 5'd6;   // 位6
        32'b00000000_00000000_00000000_001?????: code = 5'd5;   // 位5
        32'b00000000_00000000_00000000_0001????: code = 5'd4;   // 位4
        32'b00000000_00000000_00000000_00001???: code = 5'd3;   // 位3
        32'b00000000_00000000_00000000_000001??: code = 5'd2;   // 位2
        32'b00000000_00000000_00000000_0000001?: code = 5'd1;   // 位1
        32'b00000000_00000000_00000000_00000001: code = 5'd0;   // 位0
        32'b00000000_00000000_00000000_00000000: code = 5'd0;   // 位0
        default:code = 5'd0;
    endcase
end

endmodule