`timescale 1ns / 1ps

module core_top(
    input  wire        aclk,
    input  wire        aresetn,
    input  wire [ 7:0] intrpt, 
    //AXI interface 
    //read reqest
    output wire [ 3:0] arid,
    output wire [31:0] araddr,
    output wire [ 7:0] arlen,
    output wire [ 2:0] arsize,
    output wire [ 1:0] arburst,
    output wire [ 1:0] arlock,
    output wire [ 3:0] arcache,
    output wire [ 2:0] arprot,
    output wire        arvalid,
    input  wire        arready,
    //read back
    input  wire [ 3:0] rid,
    input  wire [31:0] rdata,
    input  wire [ 1:0] rresp,
    input  wire        rlast,
    input  wire        rvalid,
    output wire        rready,
    //write request
    output wire [ 3:0] awid,
    output wire [31:0] awaddr,
    output wire [ 7:0] awlen,
    output wire [ 2:0] awsize,
    output wire [ 1:0] awburst,
    output wire [ 1:0] awlock,
    output wire [ 3:0] awcache,
    output wire [ 2:0] awprot,
    output wire        awvalid,
    input  wire        awready,
    //write data
    output wire [ 3:0] wid,
    output wire [31:0] wdata,
    output wire [ 3:0] wstrb,
    output wire        wlast,
    output wire        wvalid,
    input  wire        wready,
    //write back
    input  wire [ 3:0] bid,
    input  wire [ 1:0] bresp,
    input  wire        bvalid,
    output wire        bready,

    // debug
    
    input           break_point,    //闂傚倸鍊风粈渚€骞栭锕€鐤�?柣妤€鐗忕粻楣冩煃瑜滈崜姘辨崲濞戙垹绠婚柛鎰▕閺嗐垽姊洪柅鐐茶嫰閿燂拷???闂侇剙绉寸壕濠氭煟閺冨洤浜圭€规挷绶氶弻娑㈠Ψ椤旂厧顫�???濠㈣埖鍔栭悡鐔兼煛閸愩劍绁╅柛銈嗙懇閺屾稑螣缂佹ê鍞夐梺鍝勮閸斿矂鍩ユ径濞㈢喐绗熼娑卞敳缂傚�?�鍊风欢锟犲窗閺嶎厽鐓€闁挎繂顦卞畵渚€鏌熼幑鎰靛殭缂佺姵绋掗妵鍕�?閹炬惌妫ョ紓浣虹帛閸ㄥ灝顫忛搹瑙勫枂闁告洦浜ｉ崺鍛存⒑缁嬫寧鍞夌紒顕€绠栨俊鐢稿箛椤戣姤顫嶉梺闈涚箳婵兘銆�?崨�?�樷拺闁告稑锕ゆ慨鍫㈡喐閺夊灝鏆熼柟宄邦儔�?�濡烽敂鎯у汲婵犵數鍋為崹鍫曗€﹂崶顒佸€垮瀣捣绾剧厧螞閻�?牏绠撶€殿噮鍣ｉ弻鈩冩媴鐟欏嫬纾抽梺杞扮劍閹瑰洭寮幘缁樻櫢???1闂傚倸鍊烽懗鍫曞磻閵娾晛纾块柡灞诲劜閸嬫﹢鏌�???0
    input           infor_flag,     //闂傚倸鍊风粈渚€骞栭锕€鐤�?柣妤€鐗忕粻楣冩煃瑜滈崜姘辨崲濞戙垹绠婚柛鎰▕閺嗐垽姊洪柅鐐茶嫰閿燂拷???闂侇剙绉寸壕濠氭煟閺冨洤浜圭€规挷绶氶弻娑㈠Ψ椤旂厧顫�???濠㈣埖鍔栭悡鐔兼煛閸愩劍绁╅柛銈嗙懇閺屾稑螣缂佹ê鍞夐梺鍝勮閸斿矂鍩ユ径濞㈢喐绗熼娑卞敳缂傚�?�鍊风欢锟犲窗閺嶎厽鐓€闁挎繂顦卞畵渚€鏌熼幑鎰靛殭缂佺姵绋掗妵鍕�?閹炬惌妫ョ紓浣虹帛閸ㄥ灝顫忛搹瑙勫枂闁告洦浜ｉ崺鍛存⒑缁嬫寧鍞夌紒顕€绠栨俊鐢稿箛椤戣姤顫嶉梺闈涚箳婵兘銆�?崨�?�樷拺闁告稑锕ゆ慨鍫㈡喐閺夊灝鏆熼柟宄邦儔�?�濡烽敂鎯у汲婵犵數鍋為崹鍫曗€﹂崶顒佸€垮瀣捣绾剧厧螞閻�?牏绠撶€殿噮鍣ｉ弻鈩冩媴鐟欏嫬纾抽梺杞扮劍閹瑰洭寮幘缁樻櫢???1闂傚倸鍊烽懗鍫曞磻閵娾晛纾块柡灞诲劜閸嬫﹢鏌�???0
    input  [ 4:0]   reg_num,        //闂傚倸鍊风粈渚€骞栭锕€鐤�?柣妤€鐗忕粻楣冩煃瑜滈崜姘辨崲濞戙垹绠婚柛鎰▕閺嗐垽姊洪柅鐐茶嫰閿燂拷???闂侇剙绉寸壕濠氭煟閺冨洤浜圭€规挷绶氶弻娑㈠Ψ椤旂厧顫�???濠㈣埖鍔栭悡鐔兼煛閸愩劍绁╅柛銈嗙懇閺屾稑螣缂佹ê鍞夐梺鍝勮閸斿矂鍩ユ径濞㈢喐绗熼娑卞敳缂傚�?�鍊风欢锟犲窗閺嶎厽鐓€闁挎繂顦卞畵渚€鏌熼幑鎰靛殭缂佺姵绋掗妵鍕�?閹炬惌妫ョ紓浣虹帛閸ㄥ灝顫忛搹瑙勫枂闁告洦浜ｉ崺鍛存⒑缁嬫寧鍞夌紒顕€绠栨俊鐢稿箛椤戣姤顫嶉梺闈涚箳婵兘銆�?崨�?�樷拺闁告稑锕ゆ慨鍫㈡喐閺夊灝鏆熼柟宄邦儔�?�濡烽敂鎯у汲婵犵數鍋為崹鍫曗€﹂崶顒佸€垮瀣捣绾剧厧螞閻�?牏绠撶€殿噮鍣ｉ弻鈩冩媴鐟欏嫬纾抽梺杞扮劍閹瑰洭寮幘缁樻櫢???5闂傚倸鍊烽懗鍫曞磻閵娾晛纾块柡灞诲劜閸嬫﹢鏌�???0
    output          ws_valid,       //闂傚倸鍊风粈渚€骞栭锕€鐤�?柣妤€鐗忕粻楣冩煃瑜滈崜姘辨崲濞戙垹绠婚柛鎰▕閺嗐垽姊洪柅鐐茶嫰閿燂拷???闂侇剙绉寸壕濠氭煟閺冨洤浜圭€规挷绶氶弻娑㈠Ψ椤旂厧顫�???濠㈣埖鍔栭悡鐔兼煛閸愩劍绁╅柛銈嗙懇閺屾稑螣缂佹ê鍞夐梺鍝勮閸斿矂鍩ユ径濞㈢喐绗熼娑卞敳缂傚�?�鍊风欢锟犲窗閺嶎厽鐓€闁挎繂顦卞畵渚€鏌熼幑鎰靛殭缂佺姵绋掗妵鍕�?閹炬惌妫ョ紓浣虹帛閸ㄥ灝顫忛搹瑙勫枂闁告洦浜ｉ崺鍛存⒑缁嬫寧鍞夌紒顕€绠栨俊鐢稿箛椤戣姤顫嶉梺闈涚箳婵兘銆�?崨�?�樷拺闁告稑锕ゆ慨鍫㈡喐閺夊灝鏆熼柟宄邦儔閿燂拷???
    output [31:0]   rf_rdata,       //闂傚倸鍊风粈渚€骞栭锕€鐤�?柣妤€鐗忕粻楣冩煃瑜滈崜姘辨崲濞戙垹绠婚柛鎰▕閺嗐垽姊洪柅鐐茶嫰閿燂拷???闂侇剙绉寸壕濠氭煟閺冨洤浜圭€规挷绶氶弻娑㈠Ψ椤旂厧顫�???濠㈣埖鍔栭悡鐔兼煛閸愩劍绁╅柛銈嗙懇閺屾稑螣缂佹ê鍞夐梺鍝勮閸斿矂鍩ユ径濞㈢喐绗熼娑卞敳缂傚�?�鍊风欢锟犲窗閺嶎厽鐓€闁挎繂顦卞畵渚€鏌熼幑鎰靛殭缂佺姵绋掗妵鍕�?閹炬惌妫ョ紓浣虹帛閸ㄥ灝顫忛搹瑙勫枂闁告洦浜ｉ崺鍛存⒑缁嬫寧鍞夌紒顕€绠栨俊鐢稿箛椤戣姤顫嶉梺闈涚箳婵兘銆�?崨�?�樷拺闁告稑锕ゆ慨鍫㈡喐閺夊灝鏆熼柟宄邦儔閿燂拷???

    output [31:0] debug0_wb_pc,
    output [ 3:0] debug0_wb_rf_wen,
    output [ 4:0] debug0_wb_rf_wnum,
    output [31:0] debug0_wb_rf_wdata

);
    wire rst;
    assign rst = !aresetn;

    wire icache_ren;
    wire [31:0] icache_araddr;
    wire icache_rvalid;
    wire [255:0] icache_rdata;
    wire dcache_ren;
    wire [31:0] dcache_araddr;
    wire dcache_rvalid;
    wire [31:0] dcache_rdata;
    wire [3:0] dcache_wen;
    wire [255:0] dcache_wdata;
    wire [31:0] dcache_awaddr;
    wire dcache_bvalid;

    //AXI communicate
    wire axi_ce_o;
    wire [3:0] axi_wsel;   
    //AXI read
    wire [31:0] axi_rdata;
    wire axi_rdata_valid;
    wire axi_ren;
    wire axi_rready;
    wire [31:0] axi_raddr;
    wire [7:0] axi_rlen;
    wire [255:0] dcache_axi_data_block;

    //AXI write
    wire axi_wdata_resp;
    wire axi_wen;
    wire [31:0] axi_waddr;
    wire [31:0] axi_wdata;
    wire axi_wvalid;
    wire axi_wlast;
    wire [7:0] axi_wlen;
    wire [1:0] cache_brust_type;
    assign cache_brust_type = 2'b01;   
    wire [2:0] cache_brust_size;
    assign cache_brust_size = 3'b010;

    //icache  闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??缂備胶濮甸崹鍧楀春閵忋�?�鍗抽柕蹇ョ磿閸欏棝姊虹紒妯荤閿燂�????????濠电姷顣槐鏇㈠磻閹达箑纾归柡宥庡亝閺嗘粓鏌熼悜姗嗘當缁炬儳�?遍幉鎼佹偋閸繄鐟查梺鍝勬噺閹倿寮婚妸鈺傚亞闁稿本绋戦敓锟�???闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滃繘鍩€椤掍胶鈻撻柡鍛Т閻ｅ嘲鈻庨幒瀣╂睏闂佸湱鍎ら崹鐢稿磻瀹ュ棛绡€閿燂拷?????缂佺虎鍘奸悥濂稿�??濡炪倖甯掗敃锕傛�?????闁哄洨鍋熺粔鐑樸亜閵忊€冲摵鐎规洏鍔戦�?�娆撴嚃閳哄啫顦╅梻鍌氬€搁崐椋庢濮樿泛鐒垫い鎺戝€告禒婊堟煠濞茶鐏￠柡鍛埣�?�濡烽敂鎯у箺婵＄偑鍊栭幐鍫曞垂婵犳碍鍋╅柣鎴炆戦崣蹇撯攽閻樻彃鏆為柕鍥ㄧ�??鐟欏嫭纾搁柛鏂跨Ф閹广垹鈹戠€ｎ亞顦伴梺闈涒康鐎靛苯顭囬弮鍫熲拻闁稿本鐟чˇ锔姐亜閹捐尙鐭欑€殿喖鐖煎畷褰掝敋閸涱喚绉甸梻鍌氬€烽懗鍓佹兜閸洖鐤炬繝濠傜墛閸庡孩銇勯弽顐户鐎规挷绶氶幃妤呮晲鎼粹剝鐏嶉梺鍝勬噺缁捇寮婚敓锟�?铻ｅ〒姘煎灡鍟搁梻浣告啞閻楁鎮ч悩宸綎缂備焦蓱婵绱掑☉姗嗗剰婵炲牊鍔欏娲川婵犲海鍔烽梺鍝勬媼閸嬪﹤顕ｉ锔绘晪闁�?�屽墴閻涱噣骞掗敓锟�??缁犲鏌ょ喊鍗炲闁伙絾鍎抽埞鎴︽偐缂佹ɑ閿梺绋匡攻閹倿鐛径鎰櫢闁绘ê鍟挎禍妤€鈹戦悙鏉戠仧闁搞劍妞藉畷鎰版偨閸涘﹦鍙嗗┑鐘绘涧濡繈顢撻敓锟�?闇夋繝濠傚閻帡鏌″畝瀣К缂佺姵鐩顕€鍩€椤掑倷鐒婇柨鏇炲€归悡娑㈡�?�閻愮數銆婇柛�?�尭閻ｇ兘宕堕妸锔炬殾闂備浇顕ч崙鐣�?礊閸℃稑�?堟繛鎴欏灪閺咁剟鏌ｉ弬鍨�?�闁抽攱鍨垮娲敃閵堝懍绮堕梺鍏兼た閸ㄩ亶寮查崼鏇炵鐟滃繒澹�?????闁靛鍎查崳鐑樸亜閵壯冧户缂佽鲸甯�?�畷鎺戭潩濮ｆ瑱鎷�??鐟欏嫭绀€闁靛牏枪椤曪綁骞橀钘変簻闂佺偓鑹鹃崐濠氬汲濡ゅ懏鈷掗柛灞剧懆閸忓矂寮搁鍡欑＜缂備焦锚濞搭噣鏌涢埡鍌滄创鐎规洜鍘ч埞鎴�?礃閳哄啩绨存繝鐢靛仜椤曨厽鎱ㄩ幘顕呮晞闁糕剝绋掗崑鍌炴煟閺傚灝鎮戦柣鎾寸懇濮婃椽顢橀妸褏鏆犻梺璇茬箳閿燂�??闁哄矉缍佹俊鎼佸Ω閿旇鍝楃紓鍌欐祰妞村摜鏁敓鐘茬畺闁宠桨绶￠崯鍛亜閿燂拷?閸庢娊骞冮幋锔解拻濞达絽鎲￠幆鍫ユ煟椤撶儐妲烘俊鍙夊姍�?�挳鎮㈡笟顖涚カ闂備焦瀵у濠氬�?????婵ǹ鍩栭悡娆戠磽娴ｅ顏呯┍椤栫偞鐓熼幖杈剧到閸樺瓨鎱ㄦ繝鍕笡缂佹鍠栭敓锟�?閿燂�?????濡炪倖甯掗崐鍛婄濠婂牊鐓犳繛鑼额嚙閻忥繝鏌￠崨顓犲煟鐎规洘绮忛ˇ瀵哥棯閹佸仮闁哄被鍊濋幊婵嬪级鐠恒劌甯挎俊鐐€戦崕閬嵥囬悽绋跨闁割偅娲�?崐鐑芥煟閹寸儐鐒介柛妯绘倐濮婃椽宕ㄦ繝鍌氼潎闂佸憡鏌ㄩ敓锟�???濡炪倖宸婚崑鎾剁磽�?�ュ拑韬柕鍡曠窔�?�挳濮€閳ヨ櫕鐤呴梻渚€娼ч敓锟�??缂佺姵鍨甸锝夊垂椤旇鏂€闂佸疇妫勫Λ妤呮�?�閿熺姵鍊电紒妤佺☉閹冲繘宕�?⿰鍏炬棃鏁愰崨顓熸闂佺粯鎸堕崹浠嬪蓟濞戙垹绠涢柛蹇撴憸閻╁酣姊洪崫鍕靛剱闁烩晩鍨跺濠氭晬閸曨亝鍕冮梺缁樺姦閸撴盯藝閵娧呯＝濞达綀娅ｇ敮娑㈡煟閳哄﹤鐏︽鐐插暙閳诲酣骞欓崘鈺傛珜濠电偠鎻徊浠嬪箹椤愩�?�绶ゅΔ锝呭暞閳锋帡鏌涚仦鍓ф噯闁稿繐鐭傚鎼侇敂閸涱偂绨婚梺鐟扮摠缁诲啴宕虫禒瀣厓鐟滄粓宕滃鑸靛剹??鐎规洩绻濆畷妯侯啅椤斿吋顓块梺鑽ゅТ濞诧妇绮婇弶鎳筹綁宕奸悢鍓佺畾濡炪倖鐗滈崑鐐哄极鏉堛劊浜滄い鎰╁灮瀛濋梺�?�狀潐閸ㄥ潡銆佸▎鎴犻┏閻庯綆鍋嗛弳銉╂⒒娴ｈ櫣甯涙い銊ユ噹铻炴繛鍡樻尭缁犵偤鏌曟繛鍨姉婵℃彃鐗婄换娑㈠幢濡櫣浠煎銈嗘⒐濞茬喖寮婚敐鍡樺劅闁挎繂妫欏В鍕煛鐎ｅ�?閭柟顔荤矙椤㈡稑顫濋崡鐐靛幗闂備浇顕栭崰妤呫€冮崨杈剧稏婵犻潧顑愰弫鍥煟閺傛寧鎯堥柛銈嗗笚娣囧﹪鎮�????闂佺ǹ顑呯€氼噣骞戦姀銈呯�?妞ゆ梻鍘ч悿鎯р攽閿涘嫬浜�???缂備胶绮崝妤呭焵椤掍礁鍤柛妯恒偢閹箖妫冨☉鍗炴倯闂佸憡绮堥悞锔兼嫹?閿熻棄鐭傚娲濞戞艾顣哄┑鈽嗗亝閻熝勭閹间焦鍋ㄩ柛娑橈功閸�?亶鏌ｆ惔顖滅У闁稿妫楃叅闁圭虎鍠楅悡鐔哥箾閹存繂鑸归柡�?�ㄥ€濋弻宥堫檨闁告挶鍔庣槐鐐哄幢濞戞鐛ュ┑掳鍊曢幊搴ㄦ偂閺囥垺鐓欓弶鍫ョ畺濡绢噣鏌涚€ｎ剙校缂佺粯鐩獮瀣晲閸℃瑥娑ч梺璇插閻旑剟骞�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鐗堟緲閸ㄥ倹绻濋棃娑欏窛闁绘繂鐖奸弻锟犲炊閵夈儳浠鹃梺鎶芥敱鐢繝寮诲☉姘勃闁告挆鍕珮闂佽崵濮甸崝鎺楀�?閹惰棄钃熸繛鎴欏灩缁犲鎮楅棃娑欏暈闁革綆鍠氱槐鎾寸瑹閸パ勭亶濠碘槅鍋勯崯鎾偘椤旂⒈娼ㄩ柍褜鍓熼妴浣糕枎閹炬潙娈愰梺鍐叉惈椤戝洦鎯�?繝鍥ㄢ拻闁稿本鐟х粣鏃€绻涙担鍐叉椤ゅ�?�姊绘担鍛婃儓闁瑰啿绻掗崚鎺�?箻鐠囧弶妲┑鐐村灟閸ㄥ湱绮婚敐澶嬬厽闁规澘鍚€缁ㄩ绱掗妸銉吋婵﹥妞介幃鐑芥偋閸喎鍓垫繝纰樻閸嬪懘銆冮崱娆戠焿鐎广儱顦粈鍫㈡喐韫囨洖顥氶柦妯侯棦瑜版帗鏅查柛娑卞弾濡苯鈹戦垾鍐茬骇婵＄偘绮欏濠氬焺閸愨晛顎撻梺鍛婃崄鐏忔瑩宕ョ€ｎ€棃鎮╅棃娑楃捕闂佸摜鍠愰幐鍐差嚕椤愶箑绠荤紓浣姑禍褰掓⒑閸涘﹦鎳冮柛濠傜埣�?�曟繈骞嬮敓锟�?閽冪噦鎷�??閿熷鍎遍ˇ顖涘閻樼粯鐓曢柡鍥ュ妼娴滄劙鏌涚€ｎ偅灏扮紒缁樼箓閿燂拷???闁稿绉电换娑虫�??閿熺晫枪瀛濆銈嗗灥濡繈宕哄☉銏犵闁挎梻鏅崢鍗炩攽閻樼粯娑ф俊顐ｎ殜椤㈡棃鎮介崨濠勫幍闂佸憡鍨敓锟�?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鐗堟緲閸戠姴鈹戦悩瀹犲缂佺媭鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鍓х帛閸嬫﹢鏌曢崼婵愭Ц闁绘劕锕﹂幉姝�?�?濞戞ǹ鎽曢梺鍓插亖閸庢煡鍩涢幋鐘电＝濞达絽顫栭鍛弿濠㈣埖鍔栭悡鏇㈠箹鐎涙鈽夐柍褜鍓氱换鍫ョ嵁閸愵喗鏅搁柣妯哄暱娴滄粓姊洪崗鑲┿偞闁哄懏绋栭妵鎰板礋椤栨稈鎷洪梺纭呭亹閸嬫盯宕濋敂濮愪簻闁靛闄勫畷宀嬫嫹?閿熻姤娲樺畝鎼佸箖瑜斿畷濂稿閵忊晛鏅梻鍌欑閹测剝绗熷Δ鍛偍闁绘劦鍓氬▍蹇涙⒒閸屾瑧顦﹂柟纰卞亝瀵板嫰宕堕敓锟�?閻掑灚銇勯幒鍡椾壕缂佸墽铏庨崣鍐嚕閹惰棄骞㈡繛鎴炵懅閸樻捇鎮峰⿰鍕煉鐎规洘绮撻幃銏☆槹鎼淬垺顔曞┑鐐存綑閸氬顭囧▎鎴犱笉婵炴垯鍨洪悡鏇㈢叓閸ラ鍒板ù婊勭矋缁绘稑顔忛鐓庣睄濡ょ姷鍋涢崯鎶剿�????闁哄洨鍋戦崑銏ゆ煙椤斿搫鐏╅柣锝忕節瀵墎鎷犳穱鎲嬫�??閿熻棄顫忔繝姘＜婵炲棙甯掗崢锟犳⒑缁嬫鍎嶉柛鏃€鍨甸悾鐑藉即閵忥紕鍔堕悗骞垮劚閹虫劙寮婚崼銉︾厽闁绘ê鍘栭懜顏堟煕閺傚灝顒㈢紒瀣槸椤撳吋寰勭€ｎ剙寮虫繝鐢靛█濞佳兾涢鐐嶏�?銇愰幒鎾跺帗闂備礁鐏濋鍛箔閹烘顥嗗鑸靛姈閻撱儲绻濋棃娑欘棤濠�?勬礈閹喖顫濋懜纰樻嫼闂傚�?�鐗婄粙鎺椝夊⿰鍫熺厱闁绘柨鎲＄亸锔兼嫹?閿熺瓔鍠栭�?�鐑藉极閹邦厼绶炲┑鐘插閸炴椽姊绘担铏瑰笡闁告梹顨婂顐﹀箹娴ｅ憡杈堥梺闈涚墕閹叉﹢寮�?崼鐔蜂汗闂傚倸鐗婄粙鎰柦椤忓牊鈷戦柟鑲╁仜婵�?�ジ鏌ｈ箛鏃傜疄闁诡噣绠栭幃婊堟寠婢跺瞼鏆伴梻鍌欑贰閸欏繘姊介崟顖ｆ晛闁搞儺鍓氶埛鎺懨归敐鍫綈闁稿濞€閺屾稒绻濋崘顏勨吂闁绘挶鍊栭幈銊ヮ渻鐠囪弓澹曞┑鐘殿暜缁辨洟寮拠鑼殾闁绘梻鈷堥弫宥嗘叏閿燂�??绾悂宕�?ú顏呪拻濞达絿鍎ら敓锟�??闂佸鏉垮闁瑰箍鍨归濂稿幢濞嗘ɑ绁┑鐘绘涧閸婃悂骞夐敓鐘冲亗闁哄洢鍨洪悡蹇擃熆閼哥數娲存俊缁㈠櫍閹ǹ绠涢妷鈺傤€嶉梺閫涚┒閸斿秶鎹㈠┑�?�窛妞ゆ洖鎳嶉崫妤呮⒒娴ｅ憡鍟為柣妤侇殜閹囨偐�?�割喖娈ㄩ梺鍦檸閿燂拷????婵犵數鍋炲娆擃敄閿燂拷??濮樺崬鏋庨柍瑙勫灴閺佸秹宕熼鈩冩線闂備胶枪閿曘儵宕归崹顔炬殾婵犻潧妫涢弳鍡涙煃瑜滈崜鐔肩嵁閹达箑顫呴柕鍫濇噽椤撳搫顪冮妶鍡欏缂佸鍨块敓锟�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牗顕辫閺�?喖姊荤壕瀣帯閻庤鎸烽悞锔界┍婵犲浂鏁嶆繝闈涙濮规绱掗悙顒€鍔ら柛姘儐缁岃鲸绻濋崶鑸垫櫖闂佺粯鍔曢悺銊╁汲閻樼粯鐓熼幖娣�?灱婢规﹢鏌曢崼鈶跺綊锝炶箛鏇犵＜婵☆垵顕ч鎾剁磽娴ｅ壊鍎愰悗绗涘洤纾规い鏍ㄧ〒缁犻箖鎮楀☉娆樼劷闁活厼妫涚槐鎺楊敊閻ｅ本鍣ч梺浼欑悼閸忔ê顕ｉ幘顔碱潊闁绘鏁稿澶愭⒒娴ｇǹ顥忛柛�?�噽閹广垽宕熼锝嗘櫍闂佸憡绻傜€�?囧绩娴犲鐓熸慨妤€妫楅弸娑㈡煟韫囷絼绨界紒杈ㄥ笧閹风娀骞撻幒鎾搭唲婵＄偑鍊ゆ禍婊堝疮椤栨粎鐭夐柟鐑樻煛閸嬫捇鏁愭惔婵堟晼闂佷紮绲惧钘夘潖濞差亝顥堟繛鎴炴皑閻ゅ嫰姊虹粙鍖℃敾闁绘濮撮悾鐑藉箣閿燂拷?绾惧ジ鏌ｉ幇顖氱毢妞ゆ梹鍔曢埞鎴︽�?�閸モ晝校闂佸憡鎸婚悷鈺呭箖閿燂�??椤㈡岸鍩€椤掑嫬钃熺€广儱鐗滃銊╂⒑閸涘﹥鎯堢紒鐘虫尭閻ｅ嘲饪伴崼鐔蜂簻婵犻潧鍊搁ˇ鎵礊鎼粹檧�?介柣鎰级閳绘洖霉濠婂嫮绠炵€规洘鍨块弫鎾绘偐�?�曞洤骞愬┑鐘灱濞夋盯鏁冮敓锟�??椤繈濡搁埡鍌滃幍缂備礁顑呴悘婵嬪汲閻旇櫣纾奸弶鍫涘妽鐏忔壆绱掑Δ鍐ㄦ灈鐎规洘鍎奸ˇ鎶芥煟濠垫劕娅嶆慨濠冩そ楠炴牠鎮欓幓鎺濇綂婵犵數鍋涢ˇ浼存儎椤栫儑鎷�?閿熻棄顫濋懜鍨珳婵犮垼娉涢敃銊╁箺閺囥垺鈷戦梻鍫熶緱濡插爼鏌涙惔銏犫枙妞ゃ垺鐟╅獮鍥敇閻樻鍟庨梺鍝勵槸閻楀棙鏅堕悾�?€鐭撴い鎺嶉檷娴滄粍銇勯幇鈺佺労婵�?�弶鎮傞弻宥囨嫚閼碱儷褍鈹戦鐟颁壕闂備線娼ч悧鍡椢涘畝鍕婵炲樊浜濋悡鐔兼煟濡搫甯犻柤鍓蹭邯閺屾盯寮懗顖氼伃闂佸疇顕х粔褰掔嵁閸ヮ剚鍋嬮柛顐犲灩楠炲秹姊绘担鍛婂暈闁割煈鍨跺畷鎰板冀椤愮喎浜炬慨妯煎亾閿燂拷???**********************
    wire BPU_flush;
    wire inst_rreq;
    wire [31:0] inst_addr1;
    wire [31:0] inst_addr2;
    wire [31:0] BPU_pred_addr;
    wire pi_is_exception;
    wire [6:0] pi_exception_cause; 

    wire icache_inst_valid1;
    wire icache_inst_valid2;
    wire [31:0] pred_addr1_for_buffer;
    wire [31:0] pred_addr2_for_buffer;
    wire [1:0] pred_taken_for_buffer;
    wire pi_icache_is_exception1;
    wire pi_icache_is_exception2;
    wire [6:0] pi_icache_exception_cause1;
    wire [6:0] pi_icache_exception_cause2;
    wire pc_suspend;
    wire [31:0] icache_pc1;
    wire [31:0] icache_pc2;
    wire [31:0] icache_inst1;
    wire [31:0] icache_inst2;
    //*************************************************


    // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔閹虫捇鈥�?????妞ゅ繐鎳忓畷鎶芥⒑濞茶骞栨俊顐ｇ箞瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻�???婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；婵炴垟鎳為崶顒佸仺缂佸�?�ч悗顒勬⒑閻熸澘鈷旂紒顕呭灦瀹曟垿骞囬悧鍫㈠幘缂佺偓婢樺畷顒佹櫠婵犳碍鐓曢柣鎰皺閸╋絾鎱ㄦ繝鍕笡闁瑰嘲鎳樺畷銊︾�?閸屾稒鐣肩紓鍌氬€风粈渚€骞栭銏╃劷闁炽儱纾弳锕傛煛閸ャ儱鐏╃紒鐙€鍣ｉ弻銈夊箒閹烘垵濮庨梺鍛婃尭缂嶅﹤顫忛搹瑙勫枂闁告洦鍋嗛ˇ銊╂⒑缁洘娅嗛柣妤冨Т閻ｉ攱�?�奸弶鎴犵杸闂佺粯顨呴悧蹇涘储閽樺�?介幒鎶藉磹閹版澘纾婚柟鍓х帛閻撶喐淇婇妶鍌氫壕濠碘槅鍋呯粙鎾诲礆閹烘鏁囬柕蹇曞Х椤斿﹤鈹戞幊閸婃捇鎳楅崼鏇炲偍闁归棿鐒﹂悡鐔煎箹閹碱厼鐏ｉ敓锟�??濞戙垺鐓涢柛娑卞枤缁犳绱掗鍡欑М鐎殿噮鍣ｅ畷濂告偄閸濆嫬绠伴梺璇查閸樻粓宕戦幘缁樼厓鐟滄粓宕滈悢椋庢殾濞村吋娼欓敓锟�??濡炪倖鎸炬慨瀵哥矈閿曞�?�鈷戠痪顓炴噺瑜把呯磼閻樺啿鐏╃紒顔款嚙閳藉濮€閿燂拷?閹峰姊洪崜鎻掍簽闁哥姵鎹囬崺濠囧即閻旂繝绨婚梺鍝勫€搁悘婵嬵敂椤愩倗纾奸弶鍫涘妽�?�曞矉鎷�??閿熻姤娲樼敮鎺楀煝鎼淬劌绠虫繝闈涙閺嗩參姊婚崒娆掑�??濡炪倖鍨靛Λ婵嬬嵁閹达箑鐐�???闁藉啰鍠愮换娑㈠箣濞嗗繒鍔撮梺杞扮閸熸挳寮婚敐鍛傜喓鎷犻懠顒傘偡濠电姵顔栭崰妤€煤閻斿娼栭柧蹇撴贡绾惧吋淇婇婵愬殭闂傚绉撮埞鎴︽倷閹绘帞楠囩紓渚囧枟閹瑰洭鎮伴钘夌窞闁归偊鍓欑粣娑欑節閻㈤潧孝闁哥噥鍋婂畷婵嬪川鐎涙ǚ鎷洪梻鍌氱墛缁嬪牊鎯旀搴ｇ＜闁告瑥顦伴妵婵撴�??閿熻姤娲�?崹鍧楃嵁濡吋�?�氶柤纰卞墻濡茬増淇婇悙顏庢�??閿熻棄顫忔繝姘偍鐟滄棃骞婇幘璇插�?�妞ゆ棁顫夐敓锟�??闂備礁鐤囧Λ鍕涘Δ鍛€堕柨婵嗩槹閻撳喛鎷�??閿熻棄�?�竟鍡樻櫠閺囥垺鍋傞柕鍫濐槹閻撴瑩姊婚崒姘煎殶闁告柨绉归弻宥夋煥鐎ｎ亞浼屽┑顔硷工椤嘲鐣锋總鍛婂亜闁诡厽宸婚崑鎾诲箳閹搭厾鍞甸悷婊冮鐓�???濠碉紕鏁诲畷鐔碱敍濞戞瑦鐝曢梻浣稿閻撳牓宕伴弽顐ょ�???婵﹨娅ｉ幏鐘诲灳閾忣偆浜愰梻渚婃嫹?閿熻棄鑻晶顖炴煛鐎ｎ亗鍋㈢€殿喖鎲￠幆鏃堝Ω瑜嶈ぐ鍕⒑閹肩偛鍔︽い銉︽尵缁瑦绻濆顓ㄦ嫹?閿熶粙姊婚崼鐔恒€掗柣鎺撴�?�閺屸€崇暆鐎ｎ剛蓱闂佽鍨卞Λ鍐€佸☉妯峰牚闁告稑鎷戠徊鍓ф�?????婵☆垵鍋愰悡鐘崇箾鐎涙鐭ゅù婊庝邯婵″瓨绗�?妤犵偞锚椤潡宕熼渚囨閻庤娲忛崝鎴︺€佸▎鎾崇畾鐟滃秶绮婚悙娴嬫斀闁绘ɑ顔栭弳顖涗繆閹绘帗鍤囩€规洜鎳撻悾鐑藉炊瑜嶉悘濠傤渻閵堝棛澧紒顔肩墦閹偞绻濋崶銊у弳闂佸搫娲ㄩ崑娑㈠焵閿燂�??缂嶅﹪骞冮垾鏂ユ閿燂拷?????闂備胶绮崝妤€鈻嶉妷褎鍠嗛柛鏇ㄥ墯閻濈兘姊洪崫鍕潶闁稿孩鐓￠幃鈥斥枎閹存柨浜鹃柣鐔告緲椤忣偄顭胯椤ㄥ﹤鐣烽搹顐ゎ浄閻庯綆鍋嗛崢鐢告⒑閸涘﹦鎳冩い锔藉娴滄悂鏁傞柨顖氫壕閻熸瑥瀚粈鍫ユ煕閻樺磭澧�????闂佸搫娲㈤崹鐟版纯闂傚⿴鍋勫ú锕€煤閺嶎厔鍥煛閸涱喒鎷婚梺绋挎湰閻燂妇绮婇悧鍫涗簻闁哄洤妫楅幊澶愬磻閹炬枼妲堥柟鐑樻尰閻濇艾顪冮妶鍐ㄧ仾闁荤啿鏅涢锝嗙鐎ｅ灚鏅ｉ梺缁樺姉閸庛倝鏁嶅Δ鍛拻濞达�?濮ょ涵鍫曟煕閿濆繒鐣垫鐐茬箻閿燂拷???闂備浇顕у锕傦綖婢跺⊕鍝勎熼悡搴＄亰闂佽宕�?褏绮婚弽顓熺厪閿燂�??????闂佹娊鏀遍崝娆撳蓟閻斿吋鐒介敓锟�???闁哄鍊濋弻锝夋晲婢跺瞼鏆┑顔硷功缁垶骞忛崨顖滅煓婵炲棛鍋撻ˉ鎴︽⒒娴ｅ懙褰掝敄閸涙潙绠犻幖杈剧到瀵煡姊绘担鍛婃儓缂佸绶氬畷銏ゅ箚瑜忛弳銈呫€掑锝呬壕闂佸搫鏈ú婵堢不濞戞瑧绠鹃柟顖嗗�?�顥氶梻浣藉亹閳峰牓宕滃☉銏″仼濡わ絽鍟埛鎺戙€掑锝呬壕濠电偘鍖犻崶銊ヤ罕闂佺硶鍓濈粙鎴犵不椤栫偞鐓欓悗娑欘焽缁犮儲绻涢崗鑲╁濞ｅ洤锕俊鍫曞川椤撶喐顔嶇紓浣哄亾閸庢娊濡堕幖浣歌摕闁绘梻鍘х粻鐢告煙閻戞绠撻柛鎾村▕濮婄儤�?�煎▎鎴濆煂闂佽绻戝畝鎼佺嵁閸儱惟闁挎柨澧介惁鍫ユ⒑閸涘﹤濮€闁哄�?�鍊圭粋鎺楀閵堝棌鎷洪梺闈╁瘜閸欏酣宕濆⿰鍛＜缂備焦顭囩粻鏍庨崶褝韬€规洖銈稿鎾倷閼碱剛宕洪梻鍌欑閹测剝绗熷Δ鍛；闁告洦鍨遍崐鑸点亜韫囨挻顥犵痪鎹愬亹缁辨挻鎷呯拠锛勫姺闂�?潧妫欑敮锟犲蓟閻斿壊妲归幖绮瑰椤掍降浜滈柨鏃囧Г鐏忥箓鏌″畝瀣М闁轰焦鍔欏畷銊╊敍濞嗘垿鈹忓┑锛勫亼閸婃垿宕濇繝鍥х？闁汇垻枪缁犳牗绻涢崱妯诲碍缂佺嫏鍥ㄧ厵閻庢稒顭囩粻銉︾箾閸忚偐顣插ǎ鍥э躬婵″爼宕堕‖顔哄劦閺屾冻鎷�??閿熺瓔鍋嗗ú鎾煛鐏炴枻韬柡浣瑰姈�?�板嫭绻濋崟闈涙暪婵犵數濮烽弫鍛婃叏閹绢喖鐤い鎰╁€栭浠嬫煟閹邦喖鍔嬮柛濠勬暬閺屻劌鈹戦崱娑虫嫹?閿熶粙鏌涘Ο缁樺唉閿燂�??????妞ゆ劧绲界壕鍐差渻閵堝啫鐏い銊ワ工閻ｇ兘鎮㈢喊杈ㄦ櫈闂佸吋浜介崕閬嶎敂瑜版帗鈷掑ù锝堟閸氬綊鏌涢悩鍐插闁诡喚鍏橀敓锟�????闁稿鎸搁～婵嬫偂鎼粹槅娼剧紓鍌欑贰閸犳牠鎮ч幘宕囨殾??闁糕晝鍋炲鍕传閵壯勬櫒闂傚�?�鍊风粈渚€骞栭鈷氭椽濡堕崨鍌涚☉铻栭柛娑卞弨琚濇繝纰樻閿燂�????濠碘剝褰冮悧濠囧箞閵娿儙鏃堝焵閿燂拷?铻炴繛鍡楁禋閸ゅ牊绻涘顔荤凹闁抽攱鍨垮娲敃閵堝懍绮堕梺鍏兼た閸ㄩ亶寮�????缂侇垱娲栨禍鐐箾閸繄浠㈤柡�?�⊕閵囧嫰顢橀悙鍙壭╁銈嗘穿缂嶄線鐛�?敓锟�??椤㈡瑧鍠婃潏銊хП闂傚�?�鑳堕敓锟�??濡炪倖娉﹂崶褎鐎柣鐔哥懃鐎氼喚寮�?闂備焦鐪归崹钘夘焽瑜旈崺銏ゅ醇閻旇櫣顔曟繛杈剧到閸熷潡宕㈤幑鎰╀汗闁圭儤鍨归敍婊冣攽椤曞棛鍒伴柛姘儔閹嫰顢涢悙鑼暫濠电偛妫�?ù姘跺疮閸涱喓浜滈柡鍐ㄦ处椤ュ鏌ｉ敂鐣岀煉婵﹦绮粭鐔煎焵閿燂�??椤洩顦归柟顔ㄥ洤骞㈡繛鎴烆焽閻ゅ洭姊鸿ぐ鎺戜喊闁哥姵纰嶇粙澶婎吋閸氥�?�缍婇幃鈩冩償閿濆棙鍠栭梻浣虹帛閹搁箖宕伴弽顓炶摕闁炽儱纾弳銈嗐亜閺冨洤鍚规い锔肩畱闇�???闁革綇缍�?敓锟�????闁崇粯鎹囧畷褰掝敊閻ｅ奔閭┑锛勫亼閸娿倝宕㈡ィ鍐ㄧ婵☆垯�?﹂崵鏇熴亜閹板墎鐣遍敓锟�??閸愨斂浜滈柡鍐ㄦ搐娴滃綊鏌涢弮鎾剁暠妞ゎ亜鍟存俊鍫曞幢濡ゅ啰鎳嗛梻浣告憸閸犳挻鏅跺Δ鍐焿鐎广儱顦伴敓锟�???闁�?�屽墰婢规洘绂掔€ｎ偆鍘遍柣蹇曞仦�?�曟ɑ绔熼敓锟�??閺屽秷顧�?柛鎾寸洴閿燂�????妤犵偛鍟撮幃娆撴倻濡粯鐝栭梻浣呵归張顒勫Φ濞戙垹纾婚柟鍓х帛閺呮繈鏌涚仦鐐殤闁稿﹦鍋涢�?�鍐Χ閸℃鍘愮紓浣哄У閸ㄧ數鍙呴梺鎸庢閺侇噣宕戦幘瀛樺闁告劑鍔嬪Ч妤呮⒑闁偛鑻晶顖滅磼鐎ｎ偄绗╃憸鐗堢矒濮婇缚銇愰幒鎾存殸濠碉紕鍋樼划娆忣嚕婵犳艾鐒洪柛鎰╁妿缁愮偤鏌ｈ箛鏇炰沪闁搞劍绻傞埢浠嬵敂閸涱垳鐦堥梺闈涚箞閿燂拷???婵犵妲呴崑鍛崲閸�?偞鍋╃€瑰嫭澹嬮弨浠嬫煕閿燂�??閺呮盯骞冮幋鐐电瘈闁靛骏绲剧涵鐐亜閹存繃鍠樼€规洏鍨介幃浠嬪川婵炵偓�?�奸梻浣哄帶椤洟宕愰弴銏犲嚑闁哄�?�顑欓悢鍡欐喐鎼搭煉鎷�?閿熻姤绻濋崒婊勬闂佸搫顦伴娆忣焽閵娾晜鐓曟い鎰╁€曢弸搴€亜???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鍓х帛閸嬨�?�鏌￠崘銊у闂傚偆鍨遍妵鍕即閿燂拷?娴滈箖鎮楃憴鍕闁搞劌澧庨幑銏犫攽鐎ｎ亞鍊為梺瀹犳〃閼冲爼濡堕敂鐣�?瘈缁剧増蓱椤﹪鏌涢妸褎鏆€规洘鍨块獮鍥敊绾拌鲸顥￠梻浣呵圭换妯何涚捄銊�?床闁糕剝菧娴滄粓鏌�?�鍐ㄥ闁活厼鐭傞幃浠嬵敍濞戞碍鍒涢梺鍝勮閸�?垿骞冮妶澶婄＜婵炴垶锕╅敓锟�????
    wire fb_pred_taken1;
    wire fb_pred_taken2;
    wire [31:0]fb_pc1;
    wire [31:0]fb_pc2;
    wire [31:0]fb_inst1;
    wire [31:0]fb_inst2;
    wire [1:0] fb_valid;
    wire [1:0]fb_pre_taken;
    
    
    wire [31:0]fb_pre_branch_addr1;
    wire [31:0]fb_pre_branch_addr2;
    wire [1:0] fb_is_exception1;
    wire [1:0] fb_is_exception2;
    wire [6:0] fb_pc_exception_cause1;
    wire [6:0] fb_pc_exception_cause2;
    wire [6:0] fb_instbuffer_exception_cause1;
    wire [6:0] fb_instbuffer_exception_cause2;

    wire [1:0]ex_is_bj;
    wire [31:0]ex_pc1;
    wire [31:0]ex_pc2;
    wire [1:0]ex_valid;
    wire [1:0]ex_real_taken;
    wire [31:0]ex_real_addr1;
    wire [31:0]ex_real_addr2;
    wire [31:0]ex_pred_addr1;
    wire [31:0]ex_pred_addr2;
    wire get_data_req;
    wire [7:0] flush_o;
    wire [7:0] pause_o;
    wire icacop_en;
    wire dcacop_en;
    wire [1:0]  cacop_mode;
    wire [31:0] cache_cacop_vaddr;

  
    wire  backend_dcache_ren;
    wire [3:0]  backend_dcache_wen;
    wire backend_dcache_writen;
    wire [31:0] backend_dcache_addr;
    wire [31:0] backend_dcache_write_data;

    // dcache 
    wire [31:0] dcache_backend_rdata;
    wire dcache_backend_rdata_valid;
    wire dcache_ready;

    // dcache-AXI 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�?????? cache 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栭柦鍐枛閺屾盯濡烽鐓庮潽闂佸搫鎳忛幃鍌炲蓟閵娾晜鍋嗛敓锟�??????闂傚倸鍊风粈渚€骞栭锔绘晞闁搞儺鍓欑粣妤呮煛�?�ュ骸骞栭柦鍐枛閺屻劑鎮㈤崫鍕戙垺顨ラ悙顏勭仾濞ｅ洤锕�?�娑樷攽閸℃洘鐫忛梻浣虹帛閹告悂藝闂堟侗娼栨繛宸簻娴肩�?鏌涢弴銊ュ箻濞寸厧娲娲传閵夈儛锝夋煙閸涘﹤鍔ら崡閬嶆煙閻楀牊绶茬紒鐘烘珪娣囧﹪濡堕崒姘婵＄偑鍊ら崑鍕箠閿燂拷?瀵鏁愰崨鍌滃枛閹煎綊鎯傞崫銉ь槸婵犵數鍋涢悺銊у垝閻樺磭顩查柣鎰仛椤洟鏌熼幑鎰靛殭缁炬儳鍚嬬换娑㈠幢濡桨鍒婇梺鍝ュ仜缂嶅﹤顫忛搹鍦煓婵炲棙鍎抽崜閬嶆⒑閸︻厸鎷￠柛�?�躬閻涱喛绠涘☉娆愭閿燂�?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥ｆ閺嗕即姊绘担鍛靛綊顢栭崱娑樼闁搞儺鍓欓拑鐔哥箾閹存瑥鐏╅柛妤佸▕閺屾洘绻涢崹顔煎濡炪値鍋掗崑濠傤潖濞差亜宸濆┑鐐寸閸ㄥ潡鐛�?幋锕€鐐婄憸婊冾焽閺嶎厽鐓ｉ煫鍥ㄦ尭鐢劑鏌涚€ｎ偅宕岀€规洜鍏�?、姗€鎮欓幇鍓佺М闁哄本娲熼敓锟�???闁哄棴缍�?弻鈩冩媴鐟欏嫬纾抽梺杞扮劍閹瑰洭寮幘缁樻櫢???闂傚倸鍊峰ù鍥р枖閺囥垹闂柨鏇炲€哥粻顖炴�????闂備浇顕х€涒晠顢欓弽顓炵獥闁哄稁鍘奸悿顕€鏌涜椤ㄥ懘鎮″┑瀣婵烇綆鍓欐俊鑲╃磼閻樺磭娲撮柡灞界Ф閹即鍨鹃崗鍛棜缂傚�?�鍊烽梽宥夊礉�?�€鍕舵�??閿熻棄鐣￠幏鏃€鐩畷銊╁箹椤撶喐娅囬梻渚€娼х换鍡涘焵椤掍礁澧俊鏌ヤ憾濮婄粯鎷呯粵瀣秷闂佽鍠栭崐鑽ゅ垝婵犳艾鍐€鐟滃繘寮抽敂鐣�?鐎瑰壊鍠曠花濂告煛閸涱喚鍙€闁哄本鐩崺鍕礂閿燂�??娴滄粓顢氶敐澶婄閹艰揪绲块惁鍫ユ⒑濮瑰洤鐏叉繛浣冲啰鎽ラ梻鍌欒兌閹虫捇宕捄銊�?�???闁靛棔绶氬顕€宕奸悢铚傛睏缂傚倸鍊烽悞锕傗€﹂崶顒€鍌ㄩ柣銏犳啞閳锋垿鏌ゆ慨鎰舵嫹?閿熶粙寮搁幋鐐电瘈闁靛繆妲勯懓鎸庛亜閵忊剝顥堟い銏★耿閹瑩鍩￠崒娑欐緫闂傚倷鐒﹂弸濂稿疾濞戙垹鐤い鏍仜绾惧綊鏌熼柇锕€鍘撮敓锟�??娴犲鐓ユ繛鎴灻鈺呮煕濡粯灏﹂柡灞稿墲閹峰懐绮欐惔鎾充壕闁割煈鍠氶弳锕傛煥濠靛棭妲搁崬顖炴偡濠婂啴鍙勭€殿喖寮剁缓浠嬪川婵炵偓瀚介梻浣呵归張顒勬嚌妤ｅ啫鐒垫い鎺嶇劍閸婃劧鎷�?閿熻姤娲�?崝鏍囬悧鍫熷劅闁挎繂娲ㄩ崝璺衡攽閻愬瓨灏伴柛鈺佸暣瀹曟垿骞�?幖顓燁啍闂佺粯鍔曢敓锟�???闂備浇妗ㄩ悞锕傚箲閸ヮ剙绠栭柍鍝勬噺閸ゆ垶銇勯幒鎴Ц闁轰礁缍婂濠氬磼濞嗘埈妲紓鍌氱Т閿曘�?�鐏嬮柣鐘充航閸斿酣鎯岄崱妞曞綊鏁愰崨顔兼殘缂備胶铏庨崹璺侯潖婵犳艾纾兼繛鍡樺焾濡差喚绱撻崒姘毙㈤柨鏇樺€涢悘�?�煟閻樺厖鑸柛鏂块叄閹矂宕卞鏇炵秺閺佹劙宕奸悤浣峰摋濠电偞鍨堕幐鍝ョ矓瑜版帒钃熼柍銉�?墯閸氬鏌涢幇鈺佸閹喎鈹戦悙鑼憼缂侇喖绉堕崚鎺�?箻鐠囪尪鎽曢梺璺ㄥ枔婵挳鎮欐繝鍥ㄧ厓閺夌偟澧楅ˇ閿嬬箾�?�€濠佺盎妞ゎ亜鍟存俊鍫曞礃閵娿儱袘闂備胶枪椤戝啴宕愬┑瀣祦闁告劑鍓弮鍫濈劦妞ゆ帒�?�哥紞鏍ㄧ節闂堟侗鍎愰柛濠囨敱閵囧嫰骞掗崱妞惧婵＄偑鍊曢敓锟�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴????闂傚倷绀�?幉锟犳偡閵壯勫床閿燂�???鐎殿喖顭峰鎾閻樿鏁规繝鐢靛Т閻忔岸宕濋弽銊︽珡闂傚倸鍊风粈渚€骞栭锕€绠悗锝庡亞椤╁弶銇勮箛鎾愁伌婵炲吋鐗滅槐鎾存媴閼测剝鍨堕崚濠囧箻椤旂晫鍘鹃梺璇�?�幗鐢帡宕濋妶澶嬬厪闁糕剝顨愰煬顒佹叏婵犲啯銇濇俊顐㈠暣閸╋繝宕橀顖樺€楃槐鎾存媴閸濆嫅锝夋煙閻熺増鍠橀柟顔诲嵆椤㈡瑧鎹勯妸褎婢戞繝鐢靛仦閸ㄥ爼鎮烽敓锟�??閳诲秹濮€閵堝棌鎷洪柣鐘充航閸斿苯鈻嶉幇鐗堢厵闁告垯鍊栭敓锟�????
    wire dev_rrdy_to_cache;
    wire dev_wrdy_to_cache;

    wire duncache_rvalid;
    wire [31:0] duncache_rdata;
    wire  duncache_ren;
    wire [31:0] duncache_raddr;

    wire duncache_write_finish;
    wire duncache_wen;
    wire [31:0] duncache_wdata;
    wire [31:0] duncache_waddr;
    
    wire [31:0] new_pc_from_ctrl;
    wire [1:0] BPU_pred_taken;

    //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭�??妤犵偛顦甸弫鎾绘偐閸愬弶鐤勯梻浣筋嚃閸ㄥジ鎮�?幇顖樹汗閿燂�??????缂傚倷鐒︾粙鎴︻敄閸℃稑鐤炬繝濠傚枤濞撳鏌曢崼婵囶棞缂佹甯￠幃妤€顫濋悡搴＄睄閻庤娲樺ú鏍敇閸忕厧绶為悗锝庡墮楠炲牓姊绘担鍛婅�?闁稿簺鍊楅幑銏ゅ礃閵娿垺鐏�???婵炲樊浜濋埛鎺懨归敐鍛暈闁诡垰鐗婇妵鍕晜鐠囪尙浠搁梺璇�?�暙閸曨厾鐦堥梺鎼炲�?閸滀礁鏁归梻鍌欑缂嶅﹤�??????闁诡垰鑻灃闁告侗鍠氶崢閬嶆⒑閺傘儲娅呴柛鐔跺嵆楠炲﹪宕ㄩ婊勶紡闂佽鍨庨崘鈺嬫嫹?閿熻姤绻涢敐鍛悙闁挎洦浜獮鍐ㄢ枎閹垮啯鏅㈤梺绋胯閸婃牠寮茬徊姒_addr闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏇炲€归崕鎴犳喐閻�?牆绗掗敓锟�?????闁�?�屽墴閿燂拷?閿燂�?????濡炪倖甯婄粈渚€宕甸敓锟�??闇夋繝濠傚缁犳绱掗鐣岊暡婵炵厧绻樻俊姝岊槾闁伙箑鐗撳娲箹閻愭彃濡ч梺鍛婁緱閿燂拷???闂傚倸鍊搁崐宄懊归崶褉鏋栭柡鍥ュ灩闂傤垶鏌ㄩ弴鐑囨嫹?閿熺晫绮婚鐐寸叆闁绘洖鍊归敓锟�??
    wire [31:0] csr_dmw0;//dmw0闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏃堟暜閸嬫挾绮☉妯诲櫧闁活厽鐟╅弻鐔告綇閸撗呮殸闁诲孩鑹鹃ˇ浼村Φ閸曨垰绠抽柛鈩冦仦婢规洟姊绘担鐟邦嚋婵炴彃绻樺畷瑙勭鐎ｎ亝鐎梺鐟板⒔缁垶寮查幖浣圭叆闁绘洖鍊归敓锟�??闂備浇顕х€涒晠顢欓弽顓為�???鐎规洘鍨剁换婵嬪磼濠婂嫭顔曢梻浣虹帛閹稿摜鑺遍崼鏇為唶妞ゅ繐鐗婇悡鏇熺箾閹存繂鑸归柣搴㈡そ閺屾洝绠�????闂佹娊鏀遍崹鍧楀蓟濞戞ǚ鏀介柛鈩冾殢娴犵厧顪冮妶鍛闁稿锕濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢�??27:25]闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏃堟暜閸嬫挾绮☉妯诲櫧闁活厽鐟╅弻鐔告綇妤ｅ啯顎嶉梺鎼炲€栭崝鏍Φ閸曨垰鍐€闁靛ě鍛獥濠电偛鐡ㄧ划宀€绱炴繝鍥ц摕闁挎稑�?�▽顏堟偣閸ャ劌绲诲┑顔芥礋濮婃椽骞�???????濞村吋娼欓拑鐔兼煟閺冨浄鎷�??闁稿鎸搁埥澶娾枍椤撗傜敖缂侇噮鍙€椤﹀绱掓潏銊ユ诞妤犵偛娲、妯款槼闁伙絽鐖煎濠氬炊瑜滈敓锟�?闂佸搫琚崝�?勫煘閹达箑骞㈡慨妤€妫欓敓銉╂⒒娴ｈ銇熼柛妯煎帶铻炴繝闈涱儏缁犳牜鎲搁悧鍫濈瑨缂佺姵绋掗妵鍕棘閸喗鍊梺璇茬箰閻楁捇骞冮敓锟�?閳绘捇宕归鐣屼壕闂備浇妗ㄧ粈渚€鈥�?畡鎵殾閿燂�?????濡炪倖甯婇梽宥嗙濠婂牊鐓欓柣鎴灻悘銉︺亜韫囧﹥娅婇柟顔煎槻閳诲骸鈻庨幋鐘虫婵°�?�濮烽崑鐐烘偋閺団€崇�?�婵＄偑鍊栧濠氬磻閹剧粯鐓冪憸婊堝礈濮樿埖鍋嬫繝濠傛噹閸ㄦ繂鈹戦悩鍙夌ォ闁轰礁顑夐弻宥堫檨闁告挾鍠庨锝嗙�?濮橆厼浜滈梺鍏肩ゴ閺呮稓绮婇敃鍌涒拺闁告捁灏欓崢娑㈡煕閻樺磭顣茬紒鍌涘笚缁轰粙宕ㄦ繛鐐闂備胶顢婇崑鎰板磻濞戙垹鐒甸敓锟�?????閻庤娲╃紞浣哥暦閿燂拷?閳ワ箓骞嬪┑鍥跺悪闂傚�?�绀佹竟濠囧磻閸涱劶娲�?瑜庨弳婊堟⒑閼姐倕鏋戠紒顔肩焸閺屽﹪鏁愭径濠勭暫婵°�?�绲介崯顖炴倿閿燂拷??楠炲灝鍔氭俊顐ｇ洴�?�曘垽鏌嗗鍡忔嫼闂佸湱枪鐎涒晠藟閸℃せ�?介敓锟�?????濠电偛妫庨崹钘夌暦閿濆棗绶為敓锟�???妞ゆ梹娲熷铏圭磼濡纰嶆俊銈囧У閹�?�顕ｉ幎鑺ユ櫜濠㈣泛顑囬崢闈涱渻閵堝棛澧柤褰掔畺�?�娊鏁愰崶锝呬壕閻熸瑥瀚粈鍫ユ煕閻樺磭澧甸柕鍡曠铻栧ù锝囨嚀椤庢挻淇婇悙宸剰濡ょ姴鎽滅划顓㈠焺閸愵亞鐦堥悗鍏稿嵆閺€鍗烆熆閿燂�??閿燂�??妞ゆ帊鐒︾粈瀣舵�??閿熻姤娲�?崝娆忕暦閻戠瓔鏁囬柣鏃囨閺嗐垻绱撻崒姘炬嫹?閿熶粙宕愰悜鑺ュ€块柨鏇炲€告闂佺粯鍔楅崕銈夊磹閸ф鐓ラ敓锟�?????缂備胶濯崹鍫曞蓟濞戞ǚ妲堟俊顖氬悑閹插ジ姊洪崫鍕�?櫤闁诡喖鍊垮濠氬Ω閳哄�?�浜為梺绋挎湰缁嬫垿顢�??
    wire [31:0] csr_dmw1;//dmw1闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏃堟暜閸嬫挾绮☉妯诲櫧闁活厽鐟╅弻鐔告綇閸撗呮殸闁诲孩鑹鹃ˇ浼村Φ閸曨垰绠抽柛鈩冦仦婢规洟姊绘担鐟邦嚋婵炴彃绻樺畷瑙勭鐎ｎ亝鐎梺鐟板⒔缁垶寮查幖浣圭叆闁绘洖鍊归敓锟�??闂備浇顕х€涒晠顢欓弽顓為�???鐎规洘鍨剁换婵嬪磼濠婂嫭顔曢梻浣虹帛閹稿摜鑺遍崼鏇為唶妞ゅ繐鐗婇悡鏇熺箾閹存繂鑸归柣搴㈡そ閺屾洝绠�????闂佹娊鏀遍崹鍧楀蓟濞戞ǚ鏀介柛鈩冾殢娴犵厧顪冮妶鍛闁稿锕濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢�??27:25]闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏃堟暜閸嬫挾绮☉妯诲櫧闁活厽鐟╅弻鐔告綇妤ｅ啯顎嶉梺鎼炲€栭崝鏍Φ閸曨垰鍐€闁靛ě鍛獥濠电偛鐡ㄧ划宀€绱炴繝鍥ц摕闁挎稑�?�▽顏堟偣閸ャ劌绲诲┑顔芥礋濮婃椽骞�???????濞村吋娼欓拑鐔兼煟閺冨浄鎷�??闁稿鎸搁埥澶娾枍椤撗傜敖缂侇噮鍙€椤﹀绱掓潏銊ユ诞妤犵偛娲、妯款槼闁伙絽鐖煎濠氬炊瑜滈敓锟�?闂佸搫琚崝�?勫煘閹达箑骞㈡慨妤€妫欓敓銉╂⒒娴ｈ銇熼柛妯煎帶铻炴繝闈涱儏缁犳牜鎲搁悧鍫濈瑨缂佺姵绋掗妵鍕棘閸喗鍊梺璇茬箰閻楁捇骞冮敓锟�?閳绘捇宕归鐣屼壕闂備浇妗ㄧ粈渚€鈥�?畡鎵殾閿燂�?????濡炪倖甯婇梽宥嗙濠婂牊鐓欓柣鎴灻悘銉︺亜韫囧﹥娅婇柟顔煎槻閳诲骸鈻庨幋鐘虫婵°�?�濮烽崑鐐烘偋閺団€崇�?�婵＄偑鍊栧濠氬磻閹剧粯鐓冪憸婊堝礈濮樿埖鍋嬫繝濠傛噹閸ㄦ繂鈹戦悩鍙夌ォ闁轰礁顑夐弻宥堫檨闁告挾鍠庨锝嗙�?濮橆厼浜滈梺鍏肩ゴ閺呮稓绮婇敃鍌涒拺闁告捁灏欓崢娑㈡煕閻樺磭顣茬紒鍌涘笚缁轰粙宕ㄦ繛鐐闂備胶顢婇崑鎰板磻濞戙垹鐒甸敓锟�?????閻庤娲╃紞浣哥暦閿燂拷?閳ワ箓骞嬪┑鍥跺悪闂傚�?�绀佹竟濠囧磻閸涱劶娲�?瑜庨弳婊堟⒑閼姐倕鏋戠紒顔肩焸閺屽﹪鏁愭径濠勭暫婵°�?�绲介崯顖炴倿閿燂拷??楠炲灝鍔氭俊顐ｇ洴�?�曘垽鏌嗗鍡忔嫼闂佸湱枪鐎涒晠藟閸℃せ�?介敓锟�?????濠电偛妫庨崹钘夌暦閿濆棗绶為敓锟�???妞ゆ梹娲熷铏圭磼濡纰嶆俊銈囧У閹�?�顕ｉ幎鑺ユ櫜濠㈣泛顑囬崢闈涱渻閵堝棛澧柤褰掔畺�?�娊鏁愰崶锝呬壕閻熸瑥瀚粈鍫ユ煕閻樺磭澧甸柕鍡曠铻栧ù锝囨嚀椤庢挻淇婇悙宸剰濡ょ姴鎽滅划顓㈠焺閸愵亞鐦堥悗鍏稿嵆閺€鍗烆熆閿燂�??閿燂�??妞ゆ帊鐒︾粈瀣舵�??閿熻姤娲�?崝娆忕暦閻戠瓔鏁囬柣鏃囨閺嗐垻绱撻崒姘炬嫹?閿熶粙宕愰悜鑺ュ€块柨鏇炲€告闂佺粯鍔楅崕銈夊磹閸ф鐓ラ敓锟�?????缂備胶濯崹鍫曞蓟濞戞ǚ妲堟俊顖氬悑閹插ジ姊洪崫鍕�?櫤闁诡喖鍊垮濠氬Ω閳哄�?�浜為梺绋挎湰缁嬫垿顢�??
    wire        csr_da;
    wire        csr_pg;
    wire [1:0]  csr_plv;

    //trans_addr to dcache
    wire [31:0] ret_data_paddr;
    wire [31:0] if_pred_addr1;
    wire [31:0] if_pred_addr2;

    wire icache_valid_out;

    front u_front
    (
    
        .cpu_clk(aclk),
        .cpu_rst(rst),

        .pred_taken(BPU_pred_taken),
        .pi_icache_is_exception1(pi_icache_is_exception1),     
        .pi_icache_is_exception2(pi_icache_is_exception2),
        .pi_icache_exception_cause1(pi_icache_exception_cause1),  
        .pi_icache_exception_cause2(pi_icache_exception_cause2),
        .pc_for_buffer1(icache_pc1),
        .pc_for_buffer2(icache_pc2),
        .pred_addr1_for_buffer(pred_addr1_for_buffer),
        .pred_addr2_for_buffer(pred_addr2_for_buffer),
        .pred_taken_for_buffer(pred_taken_for_buffer),
        .icache_pc_suspend(pc_suspend),
        .inst_for_buffer1(icache_inst1),
        .inst_for_buffer2(icache_inst2),
        .icache_inst_valid1(icache_inst_valid1),
        .icache_inst_valid2(icache_inst_valid2),
        .icache_valid_in(icache_valid_out),

    // *******************
        .fb_flush({flush_o[2],flush_o[0]}), //闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹瑩寮堕崹顕呭殭闂傚�?�鍊搁崐鐑芥倿閿曞�?�绠栭柛顐ｆ�?绾炬寧绻濇繝鍌滃閿燂拷?閸愨斂浜滈煫鍥ㄦ尵婢ь澁鎷�??閿熻姤娲樼划�?勫煘閹达附鏅柛鏇ㄥ亗閺夘參姊虹粙鍖℃敾闁搞劌鐏濋悾鐑藉即閵忊€虫濡炪倖甯婄粈浣规償婵犲洦鈷戦柛鎾村絻娴滄繄绱掔拠鑼㈡い顓炴喘�?�粙濡歌椤旀洟鎮楅悷鏉款棌闁哥姵娲滈懞閬嶅礂缁楄桨绨婚梺闈涱槶閸庤櫕鏅跺☉姘辩＜缂備焦顭囧ú�?�橆殽閻愬樊鍎旈柟顔界懅閹瑰嫭绗熼娑辨（婵犵绱曢崑鎴�?磹瑜忓濠冪鐎ｎ亞顔愬銈嗗姧缁犳垿鎮￠敓锟�?閺岀喐娼忛崜褏鏆犻梺缁樻惈缁绘繈寮诲☉銏犵労闁告劧缂氬▽顏嗙磽娴ｉ潧濡块柛妯犲浄鎷�?閿熶粙宕�?鍢壯囨煕閹扳晛濡兼い顒€鐗撳娲箰鎼淬垹顦╂繛�?�樼矤娴滄繃绌�????婵☆垵鍋愰幊婵嬫⒑闁偛鑻晶顔姐亜閺囶亞绉い銏�?�哺閿燂�??閿燂�???闁伙絿鍏�?幃鈩冩償濡粯鏉搁梺璇插嚱缂嶅棙绂嶅┑�?�辈妞ゅ繐鐗婇埛鎺楁煕鐏炲墽鎳呮い锔肩畵閺�?喓鍠婇崡鐐扮盎闁绘挶鍊濋弻鏇熺箾閻愵剚鐝旈梺姹囧€ら崳锝夊蓟濞戞粠妲煎銈冨妼閹虫劗鍒掓繝姘兼晬婵炴垶姘ㄩ鏇㈡倵閻熸澘顥忛柛鐘虫礈閼鸿鲸绺介崨濠勫幗闂佽宕樺▔娑㈠几濞戙垺鐓涢敓锟�?鐎ｎ剙鍩岄柧浼欑秮閺屾稑鈹戦崱妤婁患缂備焦顨忛崣鍐潖濞差亝鍋傞幖绮规濡本绻涚€涙鐭ゅù婊庝簻椤曪絿鎷犲ù瀣潔闂�?潧绻掓慨鐢杆夊┑瀣厽闁绘ê鍘栭懜顏堟煕閺傚潡鍙勭€规洘绻堥�?�娑㈡�??????婵犵數鍋涢悧鍡涙倶濠靛鍑犻柕鍫濐槸閸戠姵銇勮箛鎾跺�?闁绘挸鍟撮幃褰掑炊瑜嶇痪褔鏌涢悙宸Ш缂佽鲸甯￠幃鈺佺�???缂傚倷鑳剁划顖滄崲閸繄鏆﹂敓锟�???闁糕晪绻濆畷鎺戔槈濮橆剛顏归梻鍌氬€搁崐鎼佸磹閹间礁纾归柣鎴ｅГ閸ゅ嫰鏌涢幘鑼槮闁搞劍绻冮妵鍕�?椤愵�?绮�??濠㈣埖鍔栭悡娑㈡煕閵夈垺娅呴柛鎾讳憾閺屾盯濡堕崱妯碱槹闂佸搫鏈惄顖炪€�?弴銏℃櫜闁糕剝鐟Σ顒傜磽閸屾瑧鍔嶉柛鏃€鐗犻妴鍐幢濡皷鏀虫繝鐢靛Т濞村倿寮鍡欑闁瑰鍋熼。鏌ユ煠閸喗澶勯敓锟�?????婵☆垵鍋愰悡浣虹磽娓氬洤鏋熼柟鐟版搐椤曪絾绻濆顒€宓嗛梺鎸庣☉鐎氼噣寮堕崨濠勭瘈闁汇垽娼у瓭闂佺ǹ锕ラ幃鍌炲春濞戞瑥绶為柟閭﹀幐閹锋椽姊虹憴鍕姸濠殿喓鍊濆顐︽焼�?�ュ棛鍘遍梺鍝勫暊閸嬫捇鏌ｉ悢鍙夋珔妞ゆ洩绲剧换婵嗩潩椤撶偘绨荤紓浣哄亾婵姤銇旈幖浣哥柧閿燂拷??闁宠鍨块幃娆撳级閹寸姳妗撻梻浣藉吹閸ｃ儵宕归幏�?€浜遍梻浣告啞閸斿繘寮插┑鍫濆К闁逞屽墮閳规垿鎮欓懠顒€顣洪梺璇茬箲缁诲牆顕ｉ幖浣哥缂備焦顭囬崢閬嶆煟鎼搭垳绉甸柛�?�噹閻ｉ浠﹂悙顒€寮挎繝鐢靛Т閹冲繘顢旈悩鐢电＜閺夊牄鍔岀粭鎺楁懚閿濆鐓曢煫鍥ㄦ�?鐢爼鏌＄€ｅ墎鐣垫慨濠勭帛閹峰懘宕ㄩ棃娑氱Ш妞ゃ垺鐗犲畷鍗炩槈濡⒈鍞堕梻浣哥秺濡潡鎮為敂鍓т笉闁圭儤顨嗛埛鎺懨归敐鍛殘闁革富鍘藉畷鏌ユ煙閻楀牊绶查悷娆欑畵閹鏁愭惔婵堟晼闂佸搫妫寸粻鎾诲箖閿燂拷?閹瑩妫冨☉妤€顥氶梻浣告啞閻熴儳鎹㈤幇鏉跨厴闁硅揪闄勯崑鎰版煙缂佹ê淇�??闂備焦鐪归崺鍕垂闁�?秵鍎庢い鏍仜閽冪喖鏌ｉ弮鍫闁哄棗顑夐敓锟�???闁绘妫楅埢鎾澄旈崨顔规嫼闂佽崵鍠愭竟鍡涙晬瀹ュ鐓曢敓锟�?????婵烇絽娲ら敃顏堝箖閸ф鏁嶉柨婵嗘�?瑜斿缁樼瑹?闁�?�屽墰閸嬫盯鎳熼娑欐珷??闁哄被鍔戝鎾Ω閵堝洨娉挎俊鐐€ら崑鍕崲閹邦喖寮叉俊鐐€曠换鎰舵嫹?閿熺瓔浜炲Σ鎰板醇閺囩啿鎷洪梻鍌氱墛娓氭危閸洘鐓曢幖娣�?灮濞叉挳鏌℃担鐟板鐎规洖宕埢搴ㄥ箣椤撶偞娅楅梻鍌氬€峰ù鍥�?磻閹版澘鐓曢柛顐犲劚缁€鍫熺箾閸℃ɑ灏柛鎴犲У缁绘盯骞嬮悙鍐╁哺�?�劍绂掔€ｎ偆鍘撻梺闈涱槶閸庢娊鏁嶅澶嬬厵闁伙絽鑻埢鍫ユ煛閿燂�??閸犲酣鎮鹃敓鐘冲亱闁割偅绻冮銈夋⒒娴ｅ憡鍟為柣妤侇殜閹囨偐�?�割喖娈ㄩ梺鍦檸閸犳宕愰悜鑺モ拻闁割偆鍠嶇欢杈ㄧ箾闂傚鐭欐慨濠傤煼瀹曟帒顫濋钘変壕闁绘垼濮ら崵鍕煕閹捐尙鍔嶉柛蹇旂矒閺屾盯顢曢敐鍡欘槬??闁割偆鍠撻敓锟�?闂傚倸鐗婃笟妤呭磿閹扮増鐓曢悗锝呭閿燂�??闂佸搫琚崝鎴濐嚕閹绢喗鍊锋繛鏉戭儏娴滃墽鎲搁悧鍫濈瑨缁炬儳鐏濋埞鎴︽偐閸欏顦╅梺缁樻尰閻╊垶寮诲☉銏犵疀闁宠桨绀�?‖�?��?閿燂�??閸曨厽鍒涢梺鍝勮嫰缁夊綊寮�????妞ゅ繐妫涢幊鍡涙⒒閿燂拷?濞佳兾涘▎鎴炴殰闁圭儤顨愮紞鏍ㄧ�?闂堟侗鍎愰柡鍛�?閺屾稑鈽夐崡鐐差潻濡炪�?�鍎查懝楣冨煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁挎洏鍨归悾鐑芥偐缂佹ê浜归柣鐘叉穿閿燂�?????闂傚倷绶氶敓锟�??闂佺ǹ瀛╂竟鍡欐閺冨牆鍗抽柕蹇婃閹风粯绻涙潏鍓хК婵炲拑缍佹俊瀛樼�?閸ャ劎鍘遍梺瑙勫劤椤曨厾绮婚悙鐑樼厵妞ゆ梹鍎抽崢鎾煛娴ｇǹ鏆ｉ敓锟�??濡炪倖甯掔€氼參宕戦埡鍛厽闁硅揪绲鹃ˉ澶愭煢閸愵亜鏋涢柡灞炬礃�?�板嫬鈽夊鍡樺枠闂備礁鎲￠…鍥�?极鐠囧樊娼栨繛宸簻閹硅埖銇勯幘瀵糕姇閻庢碍鐩娲川婵炴帩浜俊鍫曞箹娴ｅ摜鐣哄┑顔姐仜閸嬫捇鏌℃担瑙勫磳闁诡喒鏅犲畷妯好圭€ｎ亙澹曢梺鍓茬厛閸嬪懘宕ｈ箛鏂剧箚妞ゆ牗绮�?敮璺好瑰⿰鍫㈢暫闁诡喗顨呴～婵嬫倷閿燂拷?閿燂�???闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹晠骞撻幒鏃戝晪闂傚�?�鍊搁崐椋庣矆娴ｈ櫣�?婂┑鐘蹭迹濞戙垹閿ら敓锟�??????闂備焦�?�уú宥夊磻閹剧粯鐓冮柦妯侯樈濡插吋銇勯敓锟�??缂嶅﹪寮�????閻庯綆鍓涢惁鍫ユ倵鐟欏嫭�?€鐎规洦鍓熼崺銉�?緞婵炪垺姊归幏鍛村川婵犲嫪澹曞┑鐘垫暩婵敻顢欓弽顓炵獥闁哄稁鍘介弲婵嬫煏婵炲灝鍔楅柡�?�Ч閺屻劌鈹戦崱妯侯槱濡炪�?�鍋呭ú鐔煎蓟閻斿吋鍊绘俊顖滃劋椤�?洟姊虹紒妯荤叆闁告艾顑夊畷鐢稿箳濡や胶鍘梺鍓插亝缁诲�?�顢楅姀銏�?�仏闁挎繂顦伴埛鎺楁煕鐏炴崘澹橀柍褜鍓涢崗姗€骞婂Δ鍛殝闁汇垹鍚€缁挳姊婚崒娆戝妽閻庣瑳鍏犻缚绠涘☉妯碱槷??闁告洦鍓欐禒濂告⒑缂佹ê鐏卞┑顔哄€濆畷鎴�?Ω閳哄倵鎷婚梺鍓插亞閸犳捇鍩ユ径鎰厽闊洦鎼煬顒佹叏婵犲啯銇濈€规洘绮撻獮鎾诲箳�?�ュ洦鏅奸梻鍌欑閹芥粍鎱ㄩ弶鎳ㄧ懓鐣￠幍铏€婚梺闈涚箞閸婃牠宕愭繝姘厱闁靛�?绲芥俊鍏笺亜???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥ｆ閺嗕即姊绘担鍛靛綊顢栭崱娑樼闁搞儺鍓欓拑鐕傛嫹?閿熷鍎遍悧婊冾瀶閵娾晜鈷戦柛娑橈攻鐏忎即鏌ｉ悢鏉戝閿燂拷?????妞ゅ繐绉电€靛矂姊洪棃娑氬婵☆偅绋掗弲鍫曟焼�?�ュ棛鍘�????閿燂�???濞寸�?浜堕弻鐔碱敊閸忓浜鹃柡鍌樺劜椤秴鈹戦绛嬫當婵☆偅鐩畷顒勬偨閸涘﹦鍘介梺缁橆焽閸庛倝濡撮崘顔藉仯闁逞屽墴閺佸啴宕掑鎲嬬吹婵犵數鍋為崹顖炲垂濞差亝鍋傞柡鍥ュ灩缁犲綊鎮�?☉娆樼劷闁宠棄顦甸敓锟�???缂侇喖鐭佽ぐ渚€姊洪幖鐐插妧鐎广儱鐗嗛幆鍫熶繆閵堝洤啸闁稿鍋ら獮鎴�?炊椤掑�?�绁﹂梺鍦劋椤ㄥ懐鐚惧澶嬬厱閿燂�??????闂佸憡姊归崹鐢革綖韫囨稒鎯為悷娆忓閻濅即姊洪悙钘夊姤婵炲懏娲熼幃妯侯吋閸滀焦�?�岄梺闈涚墕閸燁偅淇婃總鍛婄厵闁惧浚鍋撻懓鍧楁煛娴ｇ懓濮嶉柟顔界懃闇夐敓锟�????闂備浇顕ч崙鐣屽緤娴犲鍊舵慨妯挎硾閻ら箖鏌曡箛�?�舵�??閿熶粙鍩涢幋鐘电＜閻庯綆鍋勯敓锟�????闁规鍠氱壕濂告煏婵炲尅鎷�?閿熶粙鎯屽▎蹇婃�?闁斥晛鍟崐鎰版煕閳哄绡€鐎规洘甯掕灃濞达絽澹婃导鏍⒒閸屾熬鎷�?閿熺晫绮堥敓锟�?楠炲鏁嶉崟顒€搴婇梺绋挎湰婢规洟宕戦幘鎰佹僵闁绘挸娴锋禒鎼佹⒑閹稿海绠�?柛�?�ㄥ€濆顐�?礃椤旇偐锛滃┑鐐村灦閼归箖鐛�?崼銉︹拻濞达�?濮ょ涵鍫曟煕閿濆繒鐣垫鐐茬箻閿燂拷????闂傚倸鍊烽悞锕傚箖閸洖�?夐悘鐐电摂閻掍粙鏌ㄩ悢鍝勑ｉ柛�?�戦妵鍕即閿燂拷?娴滈箖鎮楃憴鍕闁挎洏鍨介妴浣糕枎閹存繃鐎抽柡澶婄墑閸斿海绮旈柆宥嗏拻闁稿本鐟х粣鏃€绻涙担鍐叉处閸嬪鏌涢埄鍐槈缂佺姷濞€閺�?喖寮堕崹顔肩导闂佹悶鍎烘禍璺何熼崟顐熸斀妞ゆ梻銆嬫Λ姘箾閸滃啰鎮奸柛鎺撳笒閳诲酣骞嬮悙鑼紡闂備線娼ц噹閻忕偠濮ら弳顖炴⒒閸屾熬鎷�??閿熺晫绮堥敓锟�?楠炲鏁�?????闂佺硶鍓濈粙鎴犵矆閸愵喗鐓ユ繝闈涙椤ョ�?鏌�???闁圭⒈鍋婇崺鐐哄箣閿旇棄浜圭紓鍌欑劍钃遍梺娆惧幖椤啴濡堕崱妤冧淮濠碘槅鍋呯换鍫濈暦閸濆嫧妲堥柕蹇曞Х椤斿﹪姊洪崷顓炰缓闁告柨鐬肩槐鐐寸節閸パ勭€梺鍦濠㈡﹢鏌嬮崶顒佺厽闁哄洦纰嶉ˇ鐑芥煕濠靛浂娈滄慨濠傛惈鏁堥柛銉戝懎濮堕梻浣规偠閸�?垶绂嶉崼鏇炵畾闁告洦鍨奸弫宥夋煟閹邦垰钄奸柟鑺ユ礋濮婃椽妫冨☉姘暫闂佺粯顨呯€氼厾绮嬪鍫涗汗闁圭儤鎸鹃崢鐢告⒑缂佹ê鐏﹂拑閬嶆煃闁垮娴柡宀嬬節瀹曢亶鍩℃担宄版瀳婵犳鍠栭敃銊モ枍閿濆绠柣妯款嚙閻忔娊鏌ц箛锝呬簽濞存粏鍩栫换婵堝枈婢跺瞼锛熼梺绋款儐椤洭宕氶幒鎴�?瀻闁规儳鍟块悗顓熶繆閵堝繒鍒伴柛鐕佸灦�?�彃鈹戠€ｎ偆鍘遍柣蹇曞仧閸嬫捇鎯冮幋鐐簻闁哄�?�灏呴煬顒佹叏婵犲啯銇濈€规洜鍏�?、姗€鎮欓弶娆炬闂傚�?�绀�?幉锟犲箰鐠囪尙鏆嗛柟闂寸閺嬩線鏌熼崜褏甯涢柡鍛�?�閺屻劑鎮ら崒娑橆伓??闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹晠骞撻幒鏃戝晪闂傚�?�鍊搁崐椋庣矆娴ｈ櫣�?婂┑鐘蹭迹濞戙垹閿ら敓锟�??????闂備焦�?�уú宥夊磻閹剧粯鐓冮柦妯侯樈濡插吋銇勯敓锟�??缂嶅﹪寮�????閻庯綆鍓涢敍鐔兼⒑闁偛鑻晶鍓х磽�?�ュ懏顥炵紒鍌氱Ч閹粓鎸婃径�?婂數闂備浇娉曢敓锟�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牓鍊楃粙蹇涙椤愩垺澶勯柟宄邦儏鐓ゆい蹇撶У閺呮粓姊洪崨濠冨闁告挻鐟х划濠囨嚋閸忓摜绠氶梺缁樺姦娴滄粓鍩€椤掍胶澧垫鐐村姈閵堬綁宕�?妸褝绱辨繝鐢靛仦閸ㄥ爼鎮烽妶鍥ㄥ床闁糕剝顭囩粻鎾呮嫹?閿熻棄澹婇崰鏇犺姳婵傚憡鐓冮梺鍨儏閻忔挳鏌￠敓锟�?閸犳牠骞婇弽顓炵厸濞达綁顥撻幑鏇炩攽閻樻鏆柍褜鍓濆▍鏇㈠磻閵夆晜鐓涢悘鐐登规晶鏌ユ煙瀹勭増鍣介柟鍙夋尦�?�曠喖顢曢悢铚傚闂佽澹嗘晶妤呮偂????闁哄洨鍋為幖鎰归悪鍛存缂佺粯鐩幃鈩冩償閿濆浂鍟嬪┑鐘殿暯閸撴繈鎮洪弴鈶哄洭骞橀鐣屽幗闂佹寧娲嶉崑鎾绘煟閿燂拷?濡繈宕洪悙鍝勭闁挎梻绮弲鈺呮⒑閸濆嫸鎷�??????缂備礁澧庨弫璇差潖濞差亜宸濆┑鐘茬箺?鐠恒劎纾奸柣妯虹－婢ь亪鏌ｉ敐鍥у幋??闂侀潧鐗嗗Λ妤佺濞差亝鈷戦柛娑橈功閳藉鎳濆畝鍕厵闁汇値鍨遍鐘电磼鏉堛劍宕岀€规洘甯掗埢搴ㄥ箣濠靛棭鐎撮梻鍌欑劍鐎笛冪暆閹间礁钃熼柨婵嗙墢閿燂拷?闂佽鍎抽悿鍥春閻愮儤鈷戦悗鍦�?�濞兼劙鏌涢妸銉�?仴闁靛棔�?�?埢搴ㄥ箻閺夋垳绮￠梺璇插缁嬫帡鏁嬮敓锟�?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牭绲鹃弲顏堟⒑閹稿海绠撴い锔跨矙�?�偊宕�?鐣屽弳闂佸搫鍟崐鐟扳枍閺囥垺鐓曢柡鍌濇硶閸╋綁鏌熼绛嬫疁闁绘侗鍣ｅ畷褰掝敊閻撳寒娼涘┑鐘殿暯濡插懘宕戦崨�?�樺仭闁靛鏅涢悡婵撴嫹?閿熷鍎遍ˇ顖烇綖閸涘瓨鐓忛柛顐ｇ箖椤ユ垿鏌熼柨�?�仢闁哄矉缍侀幃鈺呭礂閸涙澘鐒婚梻浣告啞閺屻劑鎳熼鐐茬厺鐎广儱顦粻娑㈡煟閿燂拷?閻楀繘宕㈤悽鍛娾拺闁告稑锕ら悘鐔兼煕婵犲啰澧遍柍褜鍓氶敓锟�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊炲銈嗗笒閿曪妇绮欒箛鏃傜瘈闁靛骏绲剧涵鐐亜閹存繃鍠橀柟顔炬暬瀹曞ジ寮撮悢鍝勫箞闂備焦鏋奸弲娑㈠矗閹版澘绠ｆ繝闈涘暞閻庢椽姊虹紒妯忣亪宕㈤弽顐ｅ床闁糕剝绋掗悡蹇涙煕椤愶絿绠栭柛锝嗘そ閺屾盯鏁愰崱妯镐虎闂佸搫鏈粙鎾诲焵椤掑﹦绉靛ù婊勭矒閿燂�????婵炵》鎷�??閿熺瓔鍤曞┑鐘宠壘閸楁娊鏌ｉ弮鍫缂佹劗鍋ゅ铏瑰寲閺囩偛鈷夐柦鍐憾閺岋絽鈹戦崶銊ь槹濠殿喖锕ㄥ▍锝囨閹烘嚦鐔烘嫚閸欏顔傞梻鍌欑閹芥粍鎱ㄩ悽鍛婂亱闁绘ê妯婇崵鏇炩攽閻樺磭顣查柡鍛�?�閺岋絽螣閸喚姣㈤梺鎸庣⊕缁矂鍩為幋锔藉€烽柡澶嬪灩娴犳悂姊洪幐搴㈢５闁哄懐濮撮悾鐑芥偨绾版ê浜鹃柨婵嗛�?�閺嬬喖鏌嶉柨�?�伌闁哄本绋戦埞鎴�?礋椤愩垹顫撻梻浣告惈椤戝棗螞閸愵喖钃熸繛鎴炲焹閸嬫捇鏁愰崘銊ヮ�?�闂�?€炲苯澧紒璇插€块、姘舵晲閸℃瑧鐦堝┑顔斤供閸樿棄鈻嶅⿰鍫熲拺闁告挻褰冩禍鏍煕閵娿儺鐓肩€殿喖鐖奸獮鏍ㄦ媴閸忓瀚奸梻浣告贡鏋繛鎾棑缁骞樼紒妯煎幍闂佸憡鍔樼亸娆戠不婵犳碍鐓�???婵炰匠鍥х厴闁瑰濮崑鎾绘晲鎼粹€茬爱闂佸綊�?卞钘夘潖濞差亜宸濆┑鐘插閻ｇ敻鏌ｆ惔銏犲毈闁革綇缍侀敓锟�????闁哄苯妫楅濂稿幢濞嗗繐绠為梻鍌欒兌缁垵鎽梺缁樻惈缁绘繂鐣烽敐澶婄妞ゆ牗绋撻崢闈涱渻閵堝棙纾甸柛�?�尵缁辨帡鎮╁畷鍥р拰閻庢鍣崑濠囩嵁濡偐纾兼俊顖濇〃濮规姊绘担钘変汗闁冲嘲鐗撳畷婊堟偄閸忕厧浠掗梺鐟板⒔缁垶鍩涢幒鎳ㄥ綊鏁愰崨顔兼殘闁荤姵鍔х换婵嗩嚕閹间緡鏁傞柛鈥崇箰娴滈箖鏌涢敂璇插箻闁靛棗锕弻锟犲川椤栨埃鏋呴悗瑙勬礃濡炰粙寮幘缁樺亹闁肩⒈鍓ㄧ槐鍙夌�?閻㈤潧孝闁挎洏鍊濋獮蹇ユ�??閿熺瓔鍠栭悿顕€骞栧ǎ顒€濡介柍閿嬪笒闇夐柨婵嗘噺閸熺偤鏌熼姘卞�?闁靛洤�?�伴弫鍌炲垂椤旇偐銈�?柣搴ゎ潐濞叉牜绱炴繝鍥х畺闁伙絽鐬奸惌娆撴偣閹帒濡块柡鍡╁亰濮婄粯鎷呴悜妯烘畬濡炪�?�娲﹂崣鍐ㄧ暦閹存惊鐔煎礂閻撳骸绨ラ梻浣虹�?�閸撴繆褰犳繛�?�樼矋缁捇寮婚悢鐓庣闁惧浚鍋呴悵鏃堟⒑鐠囪尙绠氶柡鍛█瀵鏁撻悩鎻掕€垮銈嗘尵婵柉鍊撮梻鍌欒兌閹虫捇宕甸弽顓炵???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鍓х帛閸嬨�?�鏌￠崘銊у缂佹劖顨婇弻鈥愁吋鎼粹€崇闂侀€炲苯澧剧紒鐘虫崌�?�濡歌閸嬫捇鏁愰崒娑欑彇缂備胶濮靛畝绋款潖妤﹁￥浜归柟鐑樻惈缁辩數绱撴担鎻掍壕婵炴挻鍩冮崑鎾绘�?????闁宠棄顦甸敓锟�?闁挎稑�?�獮鍫ユ⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ偄浜�?銈嗙墬缁海澹曟總鍛婄厪濠电偛鐏濋崝鎾煟閹惧啿鎮戦柟渚垮妽缁绘繈宕熼鐐殿偧闂備胶鎳撻崲鏌ュ箠閿燂拷?楠炲啴鎮滈挊澶岄獓闂佸壊鐓堥崯鈺呭箣閻樼數锛濋梺绋挎湰閻熴劑宕楅敓锟�??缁辨帡顢氶崨顓犱桓闂�?潧妫楅崯顖滄崲濠靛鐐婇柕澶堝灩娴滄儳霉閿濆懎顥忔繛灏栨櫊閹綊宕崟顒佸創闂佸摜鍋戦崝�?勨€旈崘顔嘉ч幖杈炬嫹?閿熻棄顫囬梻渚€娼ч悧鍡椢涢鐔侯浄闁冲搫鎳忛埛鎴︽煕韫囨挸鎮戦柕鍥ㄧ箓闇夋繝濠傛绾箖鏌ｉ敐鍥у幋妤犵偛娲、姗€鎮╅锝囦簽缂傚�?�鍊风欢锟犲磻閹烘�?堥柣鏂款殠濞兼牕鈹戦悩�?�犲缁炬儳鍚嬮幈銊ヮ潨閸℃骞嬮梺绋款儐閹瑰洭鐛弽銊�?闁告縿鍎荤槐顕€姊绘担鍝ョШ閿燂�?????濞达絽鎼ˉ姘舵煕閿旇骞愰柛瀣崌閹兘寮跺▎鍙ョ棯闂備線娼荤徊鍧椝夐幇鏉课﹂柟鐗堟緲缁犳娊鏌熺€电ǹ孝闁逞屽墰閸嬨�?�骞冨畡鎵冲牚闁告劗鍋撻埢鍫ユ�?�濞堝灝鏋熼柟顔煎€搁锝嗙鐎ｅ灚鏅ｉ梺缁樻煥閹碱偊鐛�?幇鐗堚拻濞达�?顫夐崑鐘绘煕鎼搭喖鐏︾€规洘娲熼弻鍡楊吋????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻�??閿濆骸澧伴柣锕€鐗撻幃妤冩喆閸曨剛顦ラ梺缁樼墪閸氬绌辨繝鍥ㄥ€婚柦妯猴級閵娧勫枑閿燂拷?閸曨偆鐣洪梺鎸庣箓濞层劎澹曟禒�?�厱閻忕偛澧介幊鍡樸亜閺傛妯€閿燂拷?????妞ゆ劧绲界壕鎶芥⒑閸濆嫭�?伴柣鈺婂灦閵嗕線寮撮�?鈩冩珳闂佹悶鍎滅仦鎯ф灎闂傚�?�鍊烽敓锟�????闂佺ǹ顑嗛幐鎼佹箒闂佺粯锚濡﹪宕曢幇鐗堢厽闁规儳鐡ㄧ粈�?�煙椤�?枻鑰块柟顔界懇楠炴捇骞掗崱妯虹槺濠电姵顔栭崰妤勫綘闂佸憡鏌ㄩ柊锝夌嵁婢舵劕绠瑰ù锝囨嚀娴滈亶姊洪崜鎻掍簼缂佽瀚伴幃鐑藉蓟閵夛腹鎷虹紓浣割儏閻忔繈顢楅�?掳浜滈柕濞垮劜椤ョ偟绱掑畝鍐摵缂佺粯绻堝畷鍫曗€栭顒€娲﹂悡鏇熺箾閹存繂鑸归柡�?�⊕缁绘盯宕�????濠殿喖锕ㄥ▍锝囨閹烘嚦鐔烘嫚閺屻儻鎷�?閿熻姤绻濋悽闈涗哗閻忓繑鐟╁畷浼村冀瑜滈崵鏇炩攽閻樺磭顣查柛瀣閺屾稓浠﹂崜褉妲堥敓锟�??????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵愭Т闁�?�屽墾缁犳挸鐣烽崼鏇ㄦ晢闁�?�屽墰缁鎮╃紒妯煎幈闂侀€涘嵆濞佳囧几閻斿吋鐓熼柟鎯у暱閺嗙喖鏌熼懠顒婃嫹??闂佸壊鍋呯换鍕囬鐐╂�?閿燂�????缂傚倸鐗呴敓锟�???濡炪倖宸婚崑鎾绘煕閻斿憡缍戦柣锝夋敱缁虹晫绮欏▎鐐秱闂備胶绮灙閻忓繑鐟︾粋宥嗗鐎涙ǚ鎷绘繛杈剧到閹诧繝骞嗛崼銉︾厱闁绘洑�?佹禍浼存煙椤斻劌娲ら獮銏＄箾閹寸偟鎳呴柛妯诲灴濮婃椽骞栭悙鎻掑Ф闂佸憡鎸诲畝鎼佸箖閳ユ枼妲堥柕蹇ョ磿閸�?亶姊洪棃娑辨Ф闁搞劌鎼埢宥夊川鐎涙鍘搁柣搴秵閸嬪懘藟閸儲鐓涢悘鐐插⒔閳藉鎽堕敐澶嬬叄闊洦绋堥崑鎾斥槈濮樺灈�?哄┑鐘垫暩閸庢垹寰婇挊澹濇椽濡舵径�?�珖濡炪�?�绻愰悧鍡欑不閺嶃劎绠鹃柛鈩冾殕缁傚鏌涢悢閿嬪櫤闁靛洤瀚板顕€宕掑顑跨帛濠电姰鍨婚幊鎾绘偋閸℃稑鐓�?柟�?�稿仜缁犵娀姊虹粙鍖℃敾妞ゃ劌妫濋獮鍫ュΩ閳哄倸浠虹紓浣割儓濞夋洟鎮惧ú顏呪拺缂佸瀵у﹢鐗堟叏濡ǹ濮傜€殿喗濞婇弫鍐磼濞戞艾甯鹃梻濠庡亜濞层�?�顢栭崨鏉戠劦妞ゆ帊鐒︾粈鍫㈢磼椤斿灝鍚圭紒杈ㄥ笒铻ｉ敓锟�?閹邦喚娉块梻鍌欑閹碱偊宕锕€纾归柣鐔稿閺嬪秹鏌￠崶銉ョ仾闁绘挻娲樻穱濠囶敍濠婂啫濡洪梺鍝ュ枔閸嬬喓妲愰幒鏃傜＜閿燂拷???婵犵數鍋熼崢褏鎹㈠Ο铏规殾婵犲﹤妫Σ楣冩偠濮樺墽绋诲ǎ鍥э躬閹瑩顢旈崟銊ヤ壕闁靛牆顦壕濠氭煕閺囥劌鐎柛銉ｅ妽缂嶅洭鏌曟繛褍鏈柨銈夋⒒娴ｅ摜绉烘俊顐㈡健閹偤鏁冮崒姘憋紱闂�?潧艌閺呮粓鎮￠弴鐔虹闁瑰鍎戦崗顒勬煕閺冨倸鏋涢柡灞剧☉铻ｉ柛蹇撳悑濮ｅ牆鈹戦纭锋敾婵＄偠妫勯悾鐑藉Ω閿斿墽鐦堥梺鍛婃处閸撴瑥鈻嶉幋鐐扮箚閿燂�??????闂傚倸�?�€氼厾绮╅悢鐓庡耿婵☆垳鈷堝ú鎼佹⒑瑜版帗锛熼柣鎺炵畵瀵彃饪伴崨顖滐紲濠电偞鍨堕敃鈺呭磿閹邦厹浜滈敓锟�??婵☆偄鍟～蹇涙惞閸︻厾锛滃┑鈽嗗灠閹碱偊锝炲鍛�?闁绘劖褰冮幃鎴︽煟閻�?繂鎳庨崹婵囥亜閹惧崬鐏╃紒鐘烘珪娣囧﹪濡堕崟顓炲闂佹悶鍊曢ˇ闈涱潖濞差亜浼犻柛鏇ㄥ幐閺嬪棝姊虹拠鑼闁告梹锕㈡俊鐢稿箛閺夎法顔婇梺瑙勫劤閻°劑鎮甸崘娴嬫�?闁绘﹩鍠栭悘杈ㄧ箾婢跺娲存い銏＄墵瀹曞崬鈽夊Ο鏄忕发闂備胶绮�?�鍥╁垝椤栫偛鐓曢柟杈鹃檮閻撴洘绻濋棃娑橆仼闁告梹鑹鹃湁闁绘ê纾惌�?�煏閸パ冾伃闁轰礁鍟村畷鎺戔槈濞嗘挻鏆樺┑锛勫亼閸娿�?�宕戦崟顓熷床闁圭儤姊归～鏇㈡煙閻戞ê娈鹃柣鏃傚劋鐎氭熬鎷�??閿熻棄澹婇崰鎺楀磻閹捐绠荤紓浣骨氶幏娲⒑閸涘﹦鈽夐柨鏇缁辨挸顫濋懜鐢靛幈闁瑰吋鐣崐鏍偟椤忓懌浜滈柕濠忓閹冲啴鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦�?�曞綊宕归鐐闂佸搫娲㈤崹褰掓嫅閻斿吋鐓忓璺虹墕閸斻�?�銇勯弬娆炬█婵﹥妞介獮鏍�?�閹绘帒螚闂備礁鎲℃笟妤呭窗濡ゅ拋鏁婇柡鍥╁枔閿燂拷?閻庡�?鍗抽弨鍗烆熆閿燂�??閿燂�??妞ゆ帊绀佹慨宥忔�??閿熻姤娲�?崹鍧楃嵁濡懙搴敄鐠恒劎娉垮┑锛勫亼閸婃牠宕濊�?�板﹪宕稿Δ浣稿壒闂佸湱鍎ら�?�鍡涙偂閵夆晜鐓熼敓锟�??????????濠电姷顣槐鏇㈠磻閹达箑纾归柡宓苯鏅犳繝鐢靛У閼瑰墽澹曟繝姘厵闁绘劦鍓涢弳妯好瑰⿰鍕煉闁哄矉绻濆畷鍫曞嫉閻㈠灚鏅肩紓鍌欑椤︿粙宕板Δ鍛﹂柛鏇ㄥ灠椤懘鏌嶉埡浣告殶妞わ缚鍗冲鐑樻姜閹殿噮妲梺鍝ュ枑閹稿啿鐣峰ú顏勭劦妞ゆ帊闄嶆禍婊堟煙閻戞ê鐏ラ柍褜鍓涚划顖滅矙婢跺⿴鍚嬪璺侯儑閸樼偓绻濆▓鍨灍闁告梹娲熼敓锟�??妞ゆ帊绶″▓妯侯熆鐟欏嫭�?嬮柟绋匡攻缁旂喎鈹戦崱娆懶ㄩ梺杞扮劍閸旀瑥鐣烽鍛闁革富鍘鹃埥澶娾攽閿涘嫬浜奸柛濠冩礈閹广垽骞囬鐟颁壕??闁搞儜鍐ㄦ闂備礁鎼崯鐘诲磻閹惧煄搴ㄥ炊瑜濋煬顒€鈹戦垾宕囧煟鐎规洘甯掗～婵嬵敃閵忊晜顥￠梻鍌氬€搁崐椋庣矆閿燂拷?閹潡宕堕濠勭◤婵犮垼鍩栭崝鏇㈠垂閸岀偞鐓曠憸搴ㄥΦ濠婂牆鐒垫い鎴ｆ硶椤︼箓鏌嶇拠鏌ュ弰妤犵偞锕㈤幖褰掝敃椤愶綆妫ㄩ梻鍌氬€风欢姘焽瑜旈幃褔宕卞▎灞戒壕婵鍘ч弸鐔哥箾閻撳寒鐓肩€殿噮鍣ｅ畷濂告偄閸欏顏烘繝鐢靛仩閹活亞寰婃禒瀣疅闁跨喓濮撮悿顕€鏌ｉ幇顔煎妺闁绘挻鐟х槐鎺炴�??閿熺瓔鍋掗崕銉╂煟閹剧偨鍋㈤柡宀€鍠栭�?�娆撳箚瑜嶉獮�?�⒑鏉炴壆顦﹂柛濠傛健楠炲啫鈻庨幙鍐╂櫌闂�?€炲苯澧柟顖涙⒐缁绘繈宕掑Δ浣规澑闂備胶绮崝鏍ь焽濞嗘挻鍊堕柣鏂垮悑閻撴洟鏌曟繛鍨姢缂佸妞介弻鐔碱敊閻ｅ本鍣紓浣虹帛缁诲牆鐣烽敓锟�??閺佸倻鎹勯妸褎鏅ㄩ梻鍌氬€烽懗鍫曞箠閹捐绠规い鎰╁€楅惌鎾绘煟閹达絾顥夐敓锟�?????闁�?�屽墴�?�曠喖顢楅崒姘疄濠电姵顔栭崰妤呭Φ濞戙垹纾婚柟鎹愮М閻熸壋鍫柛鈩冾焽閵嗘劕顪冮妶搴�?�簻缂佺粯鍔楅崣鍛渻閵堝懐绠伴悗姘间簽濡叉劙宕奸弴鐔叉嫼闂佸憡绋戦敃銉�?緞閸曨垱鐓曟俊顖濆吹閻帡鏌熼瑙勬珖缂佽鲸甯掕灒闁绘挸楠哥粻鐐寸節閻㈤潧啸闁轰礁鎲￠幈銊╁箻椤旇偐鏌堝銈嗙墬缁酣鎯岄崱娑欑厱闁逛即娼ч弸鐔兼煟閹惧娲撮柡灞剧☉閳藉宕￠悙鑼啋闂備胶纭堕弲顏嗗緤閸ф鐒垫い鎺嶇贰閸熷繘鏌涢悩宕囧�????闂備礁鐏濋鍕崲閸℃稒鐓熼柟杈剧到琚氶梺鍝勬噺閹倿寮婚妸鈺傚亞閿燂拷?????闂傚倸鍊风欢姘跺焵椤掑�?�浠滈柤娲诲灡閿燂拷???闁哄矉缍€缁犳盯寮崹顔芥嚈婵°�?�濮烽崑娑㈡偋閹剧繝绻嗛柟闂寸鍞銈嗘濡嫮绱撻幘缁樷拻濞达綀娅ｉ妴濠囨煕閹惧绠為柕鍡楀暣�?�曘劍娼忛崜褏鈼ゆ俊鐐€栭崝鎴�?磹濡ゅ啫顥氶柦妯侯棦瑜版帗鏅查柛娑卞弾濡苯鈹戦檱鐏忣亪锝炴径�?�攳濠电姴娲﹂崐鐑芥煙濞堝灝鏋ら柣鎾存崌閹鈻撻崹顔界亪濡炪値鍘鹃崗妯侯嚕椤愩埄鍚嬪璺猴功椤︽澘顪冮妶鍛闁瑰啿瀛╅崚濠冨鐎涙ǚ鎷洪梺鐓庮潟閸婃洖鐡繝鐢靛仩椤曟粎绮婚幒妤€桅闁圭増婢樼粈鍐┿亜閺囩偞顥犵紒�?�箻濮婃椽骞栭悙鎻掑Ф闂佸憡鎸诲畝鎼佸春濞戙垹绠ｉ柨鏃囨娴�?垶姊洪幖鐐插姷缂佸弶妞藉畷鎴�?箻缂佹ɑ鍎銈嗗姂閸婃挾鑺遍幘顔解拻闁稿本鐟ч崝宥夋煙椤旇偐鍩ｇ€规洘绻嗙粻娑㈠箻閹邦厾娲寸€规洜鍠栭、娑樷槈濡鍋呴梻鍌欒兌缁垶宕归悡骞盯宕熼敓锟�??閸旀棃姊婚崒娆戝妽閻庣瑳鍥ц摕闁靛⿵闄勫▍鐘裁归悩宸剱闁稿骸锕弻娑㈩敃閻樻彃濮曢梺鎶芥敱閸ㄥ潡寮诲☉妯锋婵鐗婇弫鐐�?閵忥絾纭鹃悗姘煎墴濠€浣糕攽閻樿宸ラ柟鍐插缁傛帟顦叉い顓℃硶閹叉挳宕熼鍌ゆЧ闁诲氦顫夐敓锟�??闁剧粯鐗曢湁闁挎繂鎳庣痪褔鎮�?顐ょ煓婵﹦绮幏鍛村川闂堟稓绉虹€殿喚鏁婚�?�妤呭礋閿燂�??娴狀參姊洪棃娴ュ牓寮插☉姘辩焼闁稿本澹曢崑鎾诲礂婢跺﹣澹曢梻浣告啞濞诧箓宕滃☉銏犲偍闁汇垹鎲￠埛鎴︽煙椤栧棗瀚々浼存⒑缁嬫鍎忛柟鍐查叄閹儳鐣￠幍顔芥畷闂侀€炲苯澧�???濡炪倖甯掗崰姘焽閹邦厾绠鹃柛娆忣檧閼板潡鏌熼鍡欑瘈闁搞劑绠栭獮鍥ㄦ媴閸涘⿴鍚欐繝鐢靛Х閺佸憡鎱ㄩ悽鍛婂殞闁诡垎鍕闂傚�?�鍊风欢姘焽瑜旇棟妞ゆ挶鍨圭壕鍧楁煙閹増顥夊ù鑲╁█楠炴牕菐閿燂拷?婵�?�粙鏌嶉柨�?�瑨闂囧鏌ㄥ┑鍡樺櫤闁哥喓鍋ら弻鐔碱敍濮樺崬鈪甸梺璇″枦濞夋盯锝炲┑瀣亗閹煎瓨绻傞弸鍫ユ煟鎼淬値娼愭繛鍙壝叅闁绘梻鍘ч拑鐔兼煕閳╁喚娈㈤柛姘儔閺屾稑鈽夐崡鐐茬闂侀€炲苯澧婚柛娆忓暙椤繘鎼归崷顓犵厯闂佸湱枪鐎涒晠骞忔潏鈺冪＝濞撴艾娲ら弸娑氱磼婢跺本鍤€闁伙綁�?辩€靛ジ寮堕幋鐘垫澑闂備胶绮�?�鍛存偋韫囨稑鍌ㄥù鐘差儐閳锋垿鎮归幁鎺戝婵炲懏鍔欓弻鐔煎礄閵堝棗顏�??闂傚倸鍊烽懗鍓佸垝椤栫儑鎷�?閿熶粙宕ㄩ鍥ㄧ☉閳藉顫濋敓锟�??閻忓﹤顪冮妶鍡樺蔼闁搞劌�?辩划濠氭惞椤愶紕绠氶梺闈涚墕鐎氼垶宕�?畝鍕厱??濞存粌鐖煎濠氭晲閸垻鏉搁梺鍝勬川閸嬫﹢宕敓锟�?椤啴濡堕崱妯垮亖闂佸憡娲︽禍鐐电不濮橆厾绡€閿燂拷?????闂佺顕滅换婵嬪箖閿熺姴�?冩い鏃囨娴�?厼鈹戦悙鍙夘棞缂佺粯鍔欓、鏃堝煛閸涱喚鍘介敓锟�????閻忓骏绠撻敓锟�???闁哥姵鐗犻妴浣糕枎閹寸偛鏋傞梺鍛婃处閸撴稖銇愰崨瀛樷拻濞达綁顥撴稉鑼磼閹绘帗鍋ョ€规洘顨呰灒闁惧繗顫夊▓楣冩⒑閸撴彃浜濇繛鍙夛耿�?�曠鎷�??閿熺瓔鍠楅悡鏇熴亜椤撶喎鐏ュù婊€绮欓弻娑㈡偄闁垮鏋犲┑顔硷工椤嘲鐣烽幒鎴僵妞ゆ垼妫勬禍鎯ь渻鐎ｎ亝鎹ｉ柣顓炴閵嗘帒顫濋敐鍛�?婵°倗濮烽崑鐐烘偋閻樹紮鎷�?閿熶粙寮撮姀鈩冩珖闂�?€炲苯澧扮紒顔碱煼閹晠鎳￠妶鍛导闂備焦鎮堕崕顖炲礉鎼淬劌鐓�?�璺虹灱绾惧ジ鏌ｅΟ铏癸紞濠�?呮暬閺岋紕浠﹂崜褉妲堥梺浼欑稻閿燂拷???濡炪倖甯掔€氼剛澹曠紒妯肩闁瑰瓨鐟ラ悘顏堟倵濮橆剚鍤囬柡宀嬬秮瀵剟宕归鏂ゆ�??閿熶粙姊虹紒妯诲蔼闁稿海鏁诲濠氭晲婢跺﹥顥濋梺鍦圭€涒晠宕曢幘缁樺€垫繛鎴炵懅缁犳绱掓潏銊ユ诞闁诡喗鐟╅�?�妤呭焵椤掑嫬绀夐柕鍫濐槹閻撴洘鎱ㄥ鍡�?⒒闁稿孩姊归〃銉╂�?�閼碱剙鈪垫繝纰樺墲閹倹淇婇柨瀣劅闁靛繆妲呭Λ鍐⒑缁洘鏉归柛�?�尭椤啴濡堕崱妤冪懆闁诲孩鍑归崣鍐ㄧ�?????妞ゅ繋鐒﹂敓锟�?闂備胶绮摫鐟滄澘鍟撮�?�鏃堝Χ婢跺鍘�???妞ゆ劧绲界喊宥咁渻閵堝骸浜濈紒璇茬墦楠炲啫鈻庨幙鍐╂櫌闂�?€炲苯澧存い銏℃閿燂拷???闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儵姊婚崒娆掑�??闂佹寧娲忛崐婵嬪灳閿燂拷?閻ｏ繝鏌囬敓锟�?濞堛劑姊虹憴鍕姸濠殿喓鍊濆鎻掆堪閸喓鍘介梺鎸庣箓閹虫劙鎮橀柆宥嗙厽??闁绘锕﹂幑銏犫攽鐎ｎ偄浠洪梻鍌氱墛閿燂�??闁靛繈鍊栭悡鏇炩攽閻樻彃鏆為敓锟�??????妞ゆ棁濮ら崐鎰攽闄囬崺鏍ь嚗閿燂�???閿濆骸澧鐐茬墛缁绘繂鈻撻崹顔界亶闂佹寧娲嶉弲鐘茬暦濠婂牊鏅濋柛灞炬皑閿涚喖妫呴銏�?�闁哄矉绲剧粋宥呪堪閸曗晙绨婚梺鍦檸閸ㄧ増鏅堕懠顒傛／妞ゆ挾鍋熼崺锝夋煛閿燂�??閸犳牠骞冮悜钘夌骇婵炲棗褰為�?顏嗙磽閸屾瑧鍔嶆い銊ョ墦瀹曚即寮�?????濠电偞鍨堕敃鈺侇焽閳哄�?�浜滈柟鍝勬娴滄儳顪冮妶鍐ㄥ姎濡ょ姵鎮傞崺鐐哄箣閿旇棄浜归梺鍓茬厛閸嬪懎袙閸曨垱鈷戠紒瀣儥閸庢劙鏌ｉ埡濠傜仸闁绘侗鍠楃换婵嬪磼濠婂嫭鐣烽梻浣告啞濞诧箓宕戦崟顖涘€垫い鎾卞灪閳锋垿鏌ら幁鎺戝壄妞ゅ繐鐓婚崶顒佸癄濠㈣埖顭囬崝鐑芥⒑閸濆嫮袪闁告柨娴风划濠氬礈瑜夐崑鎾绘偡閺夋妫岄梺鍝ュУ濞叉粓鎳為柆宥嗗殥闁靛牆鍊告禍楣冩煟閻斿搫顣奸柛鐔哄仧缁辨帞鎷犻敓锟�???閸ф鏄ラ柣鎰惈缁狅綁鏌ㄩ弮鍥棄濞存粌缍婂娲捶椤撶姴绗￠柣銏╁灡椤ㄥ懘鍩㈤幘娲绘晣闁绘鏁搁敍婊勪繆閵堝繒鍒伴柛鐕佸灦瀵啿饪伴崼鐔哄幐闂佸憡渚楅崰姘洪幘顔界厱闁冲搫鍟禒杈殽閻愬樊鍎旈柡浣稿€块幐濠冨緞閸℃ぞ澹曟俊鐐差儏缁ㄥ爼宕戦幘缁樺仭闁哄顑欏Λ�?勬⒑閸濄儱校妞ゃ劌妫濆鏌ュΨ閵夈垺鏂€闂佺粯锚閻忔岸寮抽埡鍛厱閻庯綆鍓欏暩婵炲瓨绮庢灙闁宠閰ｉ獮妯虹暦閸モ晛鐐婇梻鍌欑閹碱偆绮旈弻銉ョ閻庯綆鍓氬畷鏌ユ煕閳╁啰鈯曢柣鎾寸懅缁辨挻鎷呴棃娑氫患闂佸搫顑嗙粙鎾绘儉椤忓牆绠氱憸�?�磻閵忋�?�鐓涢敓锟�?鐎ｎ剛袦濡ょ姷鍋涘ú顓€€佸Δ鍛＜婵炴垶鐟ラ弸娑樷攽閻樺灚鏆╅柛�?�洴楠炲﹤鐣濋崟顐㈢€梺鑺ッˇ钘夘焽閺嶎厽鐓ｉ煫鍥ㄥ嚬濞兼劧鎷�?閿熻姤娲栭ˇ鐢稿蓟閺囩喓绠鹃柛顭戝枛婵洟姊虹紒妯肩細闁搞劏妫勯～蹇撁洪鍛画闂佸搫顦伴敓锟�????闂傚倷鑳堕幊鎾诲吹閺嶎厼绠�???婵犵數濮烽弫鍛婃叏閹绢喗鍎夊鑸靛姇缁狙囧箹鐎涙ɑ灏ù婊呭亾娣囧﹪濡堕崟顓炲闂佸憡鐟ョ换姗€寮婚敐澶婄闁挎繂妫Λ鍕磼閹冣挃缂侇噮鍨抽幑銏犫槈閵忕姷顓洪梺缁樺姈椤旀牠寮抽敓鐘冲€甸悷娆忓缁€鍐煟閹垮嫮绡€鐎殿喖顭烽幃銏ゅ�?????婵犵妲呴崹闈涚暦閻㈢ǹ鐭楅柛鈩冪⊕閳锋垿鏌熼懖鈺佷粶濠碉紕鏅槐鎺旀嫚閹绘帗娈诲Δ鐘靛仜閻楁挻淇婇幖浣肝ㄦい鏃囨缂傛捇姊绘担铏广€婇柛鎾寸箞閵嗗啴宕ㄩ婊€绗夐悗瑙勬礀濞层劎澹曢挊澹濆綊鏁愰崶鈺傛啒闂佹悶鍊栭悷锔界┍婵犲浂鏁冮柨婵嗘处閸掓盯姊虹化鏇熸澒闁稿鎸搁�?�鍐Χ閸℃鐟愮紓浣筋啇缁绘繂鐣烽婵堢杸婵炴垶鐟ч崢閬嶆⒑缂佹�?�鎴�?礈濮橆兘鏋旀繝濠傜墛閻撴瑦銇勯弬璇插婵炶绠撳畷鎴�?箛椤旂懓浜鹃柣鐔告緲椤ュ繘鏌涢悩鎰佹畼缂佽京鍋為幆鏃堟晲閸モ晪绱抽梻浣呵归張顒勬偡瑜斿畷婵嗩吋婢跺鐝旈梺鍛婎殘閸嬫劙寮ㄩ懞銉ｄ簻闁哄秲鍔庨埊鏇㈡�?�韫囥儳鐣甸柡宀嬬磿娴狅妇鎷犲ù�?�壕婵犻潧顑囧畵浣搞€掑锝呬壕濡ょ姷鍋炵敮锟犵嵁鐎ｎ亖鏀介柛鐘靛閸ㄥ灝顫忕紒妯肩懝闁�?�屽墮椤洩顦查摶鐐翠繆閵堝懏鍣洪柡鍛箖閵囧嫯绠涢幘鎰佷紝濠电偛鍚嬮悧妤冩崲濞戞﹩鍟呮い鏃囧吹閻╁孩绻涚壕瀣汗閿燂拷??闂佸搫鏈�?ú妯侯嚗閸曨垰閱囨繝闈涙椤ユ繈姊绘担鐟邦嚋缂佽鍊胯棟濞寸厧鐡ㄩ崑鍌炴煛閸ャ儱鐏柣鎾卞劦閺岋綁寮�?????????闂傚倸鍊峰ù鍥х暦閻㈢ǹ绐楅柛鈩冪☉绾惧潡鏌ｉ�?鈩冨仩闁逞屽厸缁€渚€锝炲┑瀣殝闁割煈鍋呴悵鍐测攽閻橆喖鐏辨繛澶嬬洴閺佸啴濡堕崶鈺冨箵濠电偞鍨堕敓锟�???闂備焦鐪归崹钘夘焽瑜嶉悺顓㈡⒑鐠囨彃顒㈤柛鎴濈秺瀹曟娊鏁愭径濠勭暰婵炴挻鍩冮崑鎿勬嫹?閿熻姤娲滈崢褔鍩為幋锕€�?冮柍鍝勫€瑰鎴濃攽閿涘嫬浜奸柛濠冪墪椤繗銇愰幒鎴濆殤缂傚倷鐒﹂�?�鍥偡鐟欏嫮绠鹃柟瀛樼懃閻忣亪鏌ｉ幘�?�樼闁哄瞼鍠栭獮鍡氼檨闁搞倗鍠愮换娑㈠箵閹烘梹鎲奸梺闈涙搐閿燂�????闂佹寧绋戠€氼參宕虫导�?�樺€甸悷娆忓閿燂�??閻庤娲﹂崜鐔煎春閵夛箑绶炲┑鐐靛亾閻庡鏌ｈ箛鏇炰沪闁稿孩濞婇、鏃堝捶椤撶姷锛濋梺绋挎湰閼归箖鍩€椤掍焦鍊愮€规洘鍔欓幃婊堟嚍????闂備焦�?�ч敓锟�????闂佸搫鎷嬫禍顏勵潖缂佹ɑ濯寸紒娑橆儏濞堫厾绱撴担铏瑰笡闁告梹娲熼幃楣冩倻缁涘鏅㈤梺鍛婃处閸嬪棝宕㈤幘顔解拺缁绢厼鎳忛敓锟�?????閿燂�??閸曨偅鐎繝鐢靛Т濞诧箓鎮￠弴鐔虹瘈闂傚牊绋掗ˉ婊勩亜韫囧鎷�?閿熶粙寮婚敓锟�??閿濆骸浜濋悘蹇ｅ弮閺屽秶鎲撮崟顐や紝閻庤娲熸禍鍫曞春閳╁啯濯撮悹鍥锋嫹?閿熻姤鍋戦梻鍌氬€搁崐椋庣矆閿燂�??楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犲閸ф绾ч柛顐ｇ濞呭洤鈽夐幘宕囆ч柡�?嬬秮閹垻绮欓幐搴ｅ浇闁荤喐绮庢晶妤冩暜濡ゅ懎鐤鹃柡灞诲劜閻撴洘绻涢幋婵嗚埞闁哄濡囬惀顏堫敇濞戞ü澹曢梻鍌氬€搁崐椋庣矆閿燂�??楠炲妾遍柟绛嬪亰濮婅櫣鎷犻垾铏亪闂佺ǹ锕ラ幃鍌炴晲閻愬墎鐤€婵炴垶鐟﹂崕顏堟⒑闂堚晛鐦滈柛姗€绠栭幃锟犲箻缂佹ǚ鎷洪梺闈╁瘜閸樻劙宕烽娑樹壕婵炴垶甯楀▍濠冾殽閻愯尙绠婚柡灞芥椤撳ジ宕辫箛鏂款伖闂傚倷绀�?敓锟�???闁诲孩绋堥弲婊冾嚗閸曨垰�?嬫い鏍ㄧ〒閸�?亶鏌ｆ惔顖滅У濞存粎鍏�?悡顒勵敆閸曨剛鍘藉┑鐐村灥�?�曨剟寮搁敂鍓х＜闁绘ê纾埥澶愭煃閽樺妲搁柍璇查叄楠炲洭顢樿閹寸兘姊婚崒姘炬嫹?閿熻棄霉閸パ€鏋栭柡鍥ュ灩闂傤垶鏌ㄩ弴鐑囨嫹?閿熺晫绮婚鐐寸叆闁绘洖鍊归敓锟�???闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩冾殔琚濋梻浣告啞閹稿爼宕濋幋锔惧祦闊洦绋掗弲鎼佹煥???闂傚倸鍊峰ù鍥р枖閺囥垹绐楃€广儱娲ら崹婵囩箾閸℃绂嬫繛鍏肩墬缁绘稑顔忛鑽ゅ嚬闂佸搫鎳忛幃鍌炲蓟閵娾晜鍋嗛柛灞剧☉閿燂拷??缂傚倸鍊搁崐椋庣矆閿燂拷?钘濋梺顒€绉撮弸渚€鎮归崶顏勭毢闁哄棴绠撻弻锟犲炊閳轰焦鐎荤紓浣稿閸嬨倝骞冨Δ鍛櫜闁告劑鍔岄�?�鍡欑磽娴ｉ潧濡兼い顓炲槻铻為柛娑欐儗閺佸啴鏌�????妞わ腹鏅犲娲偡閻�?牊鍠愰梺绋款儐閹瑰洤顕ｉ懠顒佸磯閻炴稈鍓濋～宥夋⒑闂堟盯鐛滅紒杈ㄦ礋瀹曘垺绂掔€ｎ偀鎷洪梺闈╁瘜閸樺ジ宕濈€ｎ偆绠鹃柛娆忣槺婢ь剛绱掗崒姘毙ラ柕鍥ㄥ姍楠炴帡骞樼捄鍝勭瑲闂佽崵鍠愮划宥囧垝閹惧磭鏆︽繝濠傚暊閺嬪酣鏌熺€电ǹ小缂佹顦甸幃妤呯嵁閸喖濮庡銈忓瘜閸ㄨ櫕绔熼弴銏犻敜婵°�?�鑳堕崢鍗炩攽鎺抽崐鏇㈠疮椤愶箑鐒垫い鎺戯功閸掍即鏌嶉挊澶樻Ц閾伙綁姊洪崹顕呭剳闁逞屽墮椤嘲螞閸涙惌鏁冮柕蹇婂墲閹瑩姊洪幐搴㈢８闁稿海鏁婚獮鍐ㄎ�?閻撱倖銇勮箛鎾村櫝闁归攱妞藉濠氬磼濮樺崬顤€缂備礁顑嗛幐鍓у垝婵犳碍鍊烽柣鎴烆焽閸樿鲸绻濋悽闈浶㈤柛鐔哄閺呭爼鎮介崨濠勫幈闂佸啿鎼崐璇裁虹€涙﹩娈介柣鎰▕閸庢棃鏌℃担闈╂�??閿熶粙骞冮崜褌娌柦妯侯槺閻ゅ嫭绻濋悽闈浶ラ柡浣告啞缁绘盯鍩€椤掍胶绠惧ù锝呭暱閸氭ê鈽夊Ο婊勬瀹曨亝鎷呯憴鍕彆闂傚�?�绀�?崯鍧�?箹椤愶箑绠犻煫鍥ㄧ⊕閸嬪倿鏌涢幇鍏哥凹闁哥姵鍔栫换婵囩節閸屾粌顣�???闁割偆鍠撶粻楣冩煕閳╁叐鎴犱焊娴煎瓨鐓曢悗锝庝憾閿燂�??闂佸搫鐭夌紞渚€鐛敓锟�??閹煎綊顢曢敐鍛存７闂傚�?�绀�?幖顐⑽涚€靛摜涓嶉柟鎹愵嚙閽冪喖鏌ｉ弬鍨�?�闁稿顑夐弻娑㈩敃閵堝懏鐏�?梺鍛婂煀缁绘繂顫忛搹瑙勫磯闁靛ǹ鍎查悵銏ゆ⒑閻熸澘娈�???闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗ù锝呮贡閻濊泛鈹戦悩鍙夊闁稿鍊块弻娑㈩敃閻樻彃濮庣紒鐐�?劤椤兘寮诲☉銏犲嵆闁靛ǹ鍎虫导鍥⒑鏉炴壆顦﹂柛濠傛健�?�濡搁埡鍌氫簽闂佺ǹ鏈敓锟�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨圭粻璇裁归敐鍫綈闁靛洦绻冮妵鍕閳╁喚妫冮悗瑙勬磸閸�?垿銆佸Ο琛℃斀闁割偆鍠愬В搴ㄦ⒒閸屾熬鎷�??閿熶粙宕愭搴ｇ�???妤犵偞鐗犻�?�鏇氱秴闁搞儺鍓欑粻銉︺亜閺冨�?�鍤€濞存粌澧界槐鎺懳旀担琛℃闂佺ǹ锕ら…宄邦嚕娴兼潙纾奸柣鎰ˉ閹峰姊虹粙鎸庢拱闁煎綊绠栭敓锟�??妞ゆ帒鍊搁崢鎾煙椤�?儳浠遍柡浣稿暣�?�曟帒顫濇潏鈺傛瘒闂傚�?�绀佹竟濠囧磻閸涱劶娲�?椤撶偛鐎梺绋挎湰椤曢亶寮崼鐔告珖婵炴挻鑹鹃敃顏堟偘濠婂嫮绠鹃悗娑欘焽閻﹦绱撳鍜冭含鐎殿喛顕ч埥澶愬閻樼數鏉搁梻鍌氬€搁悧濠勭矙閹烘鍊剁€广儱顦伴埛鎴犵磼鐎ｎ偒鍎ラ柛搴＄焸閺岋繝宕ㄩ鐐�?????婵﹥妞介獮鎰償閿濆洨鏆ら梻浣烘嚀閸熷潡鏌婇敐鍜佸殨闁规儼濮ら崑鍕煕韫囨艾浜归柛妯圭矙濮婃椽妫冨☉姘暫闂佺ǹ锕ら幉锛勭矉瀹ュ绠氱憸澶愬绩娴犲鐓熸俊顖濇娴犳盯鏌￠崱蹇旀珚閿燂拷?????閿燂�???閿燂�??????闁哄洨鍋熺粔鐚存�??閿熻姤娲栭妶绋款嚕閹绢喗鍋勯柧姘�?€婚弫楣冩⒒閸屾瑧鍔嶉悗绗涘厾娲冀椤撶偟锛欓梺鍛婄缚閸庨亶藟濮樿埖鐓欑紒�?�硶閺勫�?�霉濠婂嫮鐭掗柣鎿冨亰�?�曞爼濡搁敓锟�?闂夊秹姊洪棃鈺冨埌闁硅姤绮庡Σ鎰板箳閿燂拷?鐎氭岸鏌涘▎蹇ｆ▓婵☆偓绠撳娲传閸曨剚鎷卞┑鐐跺皺閸犲酣鎮鹃悜鑺ュ亗閹煎瓨蓱閿燂�??闂備礁澹婇崑渚€宕洪崟顖氳埞婵炲樊浜濋埛鎺懨归敐鍛暈闁哥喓鍋ら幃浠嬵敍濮樻崘鍚悗瑙勬穿缁绘繈鐛惔銊�?癄濠㈣泛瀛╅幉鐗堢節閻㈤潧浠﹂柛顭戝灦�?�曠懓煤椤忓嫮锛涢梺绯曞墲椤﹂缚銇愰幒鎾存珳闂佸憡渚楅崰妤呭窗閹邦厾绠鹃悗鐢登规牎闂佽鍠栭崐鍧楃嵁閸愩剮鏃堝焵椤掑嫬鐓濋柟鎹愵嚙閸ㄥ�?�銇勯弮鍌涙珪濞存粌鐖煎缁樻媴閾忕懓绗￠梺鐟版啞閹告娊宕�?濡炪倖宸婚崑鎾剁棯缂併垹寮€殿喗濞婇弫鍌涙叏閹邦亞鐩庨梻浣筋潐濠㈡ɑ鏅舵惔銊�?仼闂侇剙绉撮懜瑙勩亜閺嶎偄浠﹂柛瀣у墲缁绘繃绻濋崒姘缂備胶濮撮…鐑藉蓟閳╁啯濯撮柛婵勫剾閵忊槅娈版い蹇撳暙瀹撳棴鎷�??閿熻姤娲栭妶鎼佸箖閵忋�?�鐭�?璺衡看娴兼牠姊婚崒姘炬�??閿熺晫绮堥敓锟�?楠炲鏁嶉崟顓犵厯闂佺鎻梽鍕疾濠靛鐓ラ敓锟�?????缂備胶濮烽敓锟�?闁哄本鐩獮鍥Ω閿旇姤绶┑鐐茬摠缁秶鍒掗幘璇茶摕闁靛ň鏅涚猾宥夋煕閵夈劍纭炬繛鍫弮濮婅櫣鎷犻懠顒傜杽闂佺ǹ娴烽弫璇差嚕鐠囧樊鍚嬪鑸瞪戦弲婊堟⒑缁洖澧查柣鐔村€濋幖鐟邦啅濮婃瑩姊婚崒姘炬嫹?閿熶粙宕愰幖浣哥９闁归棿�?佺壕褰掓煙闂傚顦︾痪鎯х秺閺�?喖姊荤€靛壊妲紒鐐�?劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻�??閿濆骸澧伴柣锕€鐗撻幃妤冩喆閸曨剛顦ラ梺缁樼墪閸氬绌辨繝鍥ㄥ€婚柦妯猴級閵娧勫枑閿燂拷?閸曨偆鐣洪梺鎸庣箓濞层劎澹曟禒�?�厱閻忕偛澧介幊鍡樸亜閺傛妯€閿燂拷?????妞ゆ劧绲界壕鎶芥⒑閸濆嫭�?伴柣鈺婂灦閵嗕線寮撮�?鈩冩珳闂佹悶鍎滅仦鎯ф灎闂傚�?�鍊烽敓锟�????闂佺ǹ顑嗛幐鎼佹箒闂佺粯锚濡﹪宕曢幇鐗堢厽闁规儳鐡ㄧ粈�?�煙椤�?枻鑰块柟顔界懇楠炴捇骞掗崱妯虹槺濠电姵顔栭崰妤勫綘闂佸憡鏌ㄩ柊锝夌嵁婢舵劕绠瑰ù锝囨嚀娴滈亶姊洪崜鎻掍簼缂佽瀚伴幃鐑藉蓟閵夛腹鎷虹紓浣割儏閻忔繈顢楅�?掳浜滈柕濞垮劜椤ョ偟绱掑畝鍐摵缂佺粯绻堝畷鍫曗€栭顒€娲﹂悡鏇㈡倶閻愭彃鈷旈柣鎿冨灠椤法鎲撮崟顒傤槰婵烇絽娲ら敃顏堝箖濞嗘搩鏁傞柛鏇樺妼娴滈箖鏌曢崼婵囶棤妞も晛寮剁换婵囩�?閸屾粌顣洪梺姹囧€ら崰鏍箒闂佺ǹ绻愰崥�?�礊閹达附鐓熼柟鐑樺灩娴犳盯鏌曢崶褍顏鐐村浮楠炲顢涘顒夋浆缂傚倸鍊风粈渚€藝闂堟侗鐒界憸鏂匡�?�娴ｇ硶�?介柣妯款嚋�?�搞儵鎮�?鐓庢珝闁诡垰鐭傞獮鎺懳�?担鍝勫箥婵＄偑鍊栭悧妤呮偡瑜忕划锝夊棘鎼存挻鏂€闂佹枼鏅涢崯顖炲磹閹扮増鐓曢柍鍝勵儑閿燂�??閻庤娲�?敓锟�???闂佸憡鍔戦崝搴敊閸ヮ剚鈷掗柛灞捐壘?閻戣姤鍤勯柛鎾茬劍閸忔粓鏌涢锝嗙閿燂�??閸喓绡€闂傚牊渚楅崕宀勬煃瑜滈崜銊х不閹惧磭鏆﹂柛顐ｆ处閺佸棗霉閿濆毥瑙勭珶閹烘鈷掑ù锝呮啞鐠愶繝鏌涙惔娑虫�??閿熶粙濡撮崘顔煎耿婵炴垶鐟ユ禍妤€鈹戦悙鏉戠仧闁搞劍妞藉鏌ュ箹娴ｅ湱鍙嗛梺缁樻�?閿燂�?????闂傚倸鍊风欢姘跺焵椤掑�?�浠滈柤娲诲灡閺呰鎷�?閿熺晫纭堕崑鎾舵喆閸曨剛锛涢梺鍛婎殕婵炲﹪鎮伴敓锟�?閿燂�????閿燂�??閸屾稏浜滈柟鎵虫櫅閻忣亪鏌涢悩绛硅€块柡�?€鍠栭�?�娆撳Ω閵夛附鎮欓梻浣稿船濞差參寮婚敐澶婃闁割煈鍠椾簺濠电姷顣介崜婵囩箾婵犲偆娼栫紓浣股戞刊鎾煕濠靛棗顏х紓鍌涙崌濮婅櫣绮欓崸妤€寮版繛瀛樼矎濞夋盯鎮鹃悜绛嬫晬婵犲﹤�?�壕顖炴⒑闂堟丹娑㈠磼濠婂懏鍠掗梻鍌氬€烽悞锔兼嫹?閿熺獤鍛床闁稿瞼鍊涢崶銊ヮ嚤闁哄鍨归崢閬嶆⒑閸︻厼鍔嬮柛銈嗕亢閵囨劙骞掗幘�?�樼彸闂備礁澹婇崑鍛垝閹惰棄绠荤紓浣诡焽閸橆亪姊虹化鏇炲⒉妞ゃ劌鎳樺鎶芥晲婢跺鍘�??閻庯綆鍓涜ⅵ婵°�?�濮烽崑鐐垫暜閿熺姴绠栨繛鍡樻尰閸嬨劑鏌涢�?�鎴濅簼妞ゆ梹鎸搁埞鎴炲箠闁稿﹥顨嗛幈銊╂�?�閽樺锛涢梺缁樺姇閹碱偊宕归崒鐐寸厱妞ゎ厽鍨甸弸銈夋煛閸☆厾鐣甸柡�?€鍠栭�?�娑㈡�?�闊厼鏋堟繝纰夋嫹?閿熻棄�?�庨柛鏃€鍨甸～蹇撁洪鍕啇闂佺粯鍔栫粊鎾磻閹捐鍐€妞ゎ剨鎷�?閿熻姤鎯堟い顐ｇ矒閿燂拷?妞ゆ帊妞掔换鍡涙煟閵忊懚鍦矆鐎ｎ偁浜滈柡宥冨妽閻ㄦ垶銇勯弬鍖¤含婵﹥妞介幃鐑藉箥椤旇姤鍠栫紓鍌欐祰椤曆呯矓閻㈢數鐭夐柟鐑樻尵闂勫嫰鏌涘☉姗堝姛闁告﹢浜跺娲濞戣鲸顎嗛梻鍌氬鐎氼喗绂嶉幖浣规櫆闁兼亽鍎卞鎸庣節閻㈤潧孝闁瑰啿绻�?、鏃堟偐缂佹鍘遍梺鍝勭Р閸斿孩鏅�?????妞ゆ棁濮ょ亸锕傛煙椤旂晫鎳冮敓锟�?????妞ゆ劑鍨昏ぐ鎯�?攽閻樻鏆滅紒杈ㄦ礋瀹曟垿骞嬮敓锟�?绾惧綊鏌�????閿燂�??????闁�?�屽墴閿燂拷?妞ゆ帒�?�粻鏌ユ煏韫囧鎷�??閿熺晫绮婚敐鍡愪簻闁哄秲鍔庨埥澶嬨亜????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牗顕辫閺�?喖姊荤壕瀣帯閻庤鎸烽悞锔界┍婵犲浂鏁嶆繝闈涙濮规绱掗悙顒€鍔ら柛姘儐缁岃鲸绻濋崶鑸垫櫖闂佺粯鍔曢悺銊╁汲閻樼粯鐓熼幖鎼線娴溿垺淇婇銏狀伃闁糕晝鍋ら獮�?��?????闂備礁鍚嬮幃鍌氼焽瑜嶉埥澶庮樄婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閸ゆ牠骞�???婵犵數濮烽弫鍛婃叏閻㈠壊鏁婇柡宥庡幖缁愭鏌熼幑鎰靛殭缁炬崘顫夋穱濠囧Χ閸屾矮澹曢梻浣哥枃濡嫰藝閻㈢ǹ绠栭柣锝呯灱閻瑩鏌涜椤ㄥ懘寮ぐ鎺撯拻濞达絽鎲￠幆鍫熺箾鐏炲倸濮傜€规洑鍗抽獮妯兼嫚閹绘帒浜堕梻鍌欑贰閸撴瑧绮旈悽绋跨厱闁瑰濮风壕钘壝归敐鍛暛闁逞屽墯鐢繝骞冮悜钘夌閿燂�??????闂傚倷绀�?幖顐⒚洪妸鈺佺；闁绘梻鍘уЧ鏌ユ煥閺囩儑鎷�?閿熶粙鎮￠妷鈺傜厽闁哄洨鍋�???????闂傚倸鍊风欢姘跺焵椤掑�?�浠滈柤娲诲灡閺呭爼宕ｆ径鍫滅盎濡炪倖鍔戦崺鍕ｉ幖浣瑰亗闁靛牆顦伴悡鍐煕濠靛棗顏╅敓锟�?????闁哄洨鍋涚痪褏绱掔紒妯肩疄婵☆偄鍟埥澶愬础閻愭彃顥愰梺璇叉唉椤骞愭搴㈩偨婵ê澧庡畵渚€鏌″搴ｄ粓閹兼惌鐓堥弫鍡涙煃瑜滈崜姘┍婵犲啰顩烽悗锝庡亞閸�?亶姊洪棃娑氬闁硅櫕鍔栭弲銉╂⒒娴ｅ憡鎯堥柡鍫墮鐓ゆ俊顖欒閸ゆ鏌涢弴銊ヤ簮婵℃彃鐗撻弻鏇＄�?婵犲喚娼戦敓锟�????缂佸鎳撻～蹇涙惞閸︻厾锛滃┑鈽嗗灥閸嬫劙鎮鹃悜妯肩瘈闁汇垽娼ф禒婊堟煥閺囨﹫鎷�?閿熶粙鏁愰悙鍓佺杸闁哄洨濮烽敍婊冣攽閳藉棗鐏ラ柛瀣姍閹線宕奸妷锔惧幍闂佸吋绁撮弲鐐舵＂闂備緤鎷�?閿熻棄鑻晶鏌ユ倶韫囨梻鎳囬柟顖氬閹棃濮€閵忋垻妲囬梻浣圭湽閸ㄨ棄顭囪缁傛帡鍩￠崒妯圭盎闂佸搫娲ㄩ崰鎾绘儗閿燂�??缁辨帡顢欑喊杈╁悑濡ょ姷鍋為敃銏ょ嵁閸ャ劍濯撮柛娑樷看閸氭瑦绻濋悽闈浶ラ柡浣告啞閹便劑鎮介崨濠傛疄闂佺粯鍔﹂崜娆撳礉閺冨牊鈷掗柛灞剧懅椤︼箓鏌涢悢閿嬪仴妤犵偞鐗犻�?�鏇㈡晜閼恒儲鐝栭梻渚€娼чˇ顐�?疾濞戙垺鍋柣鎰靛墰閿燂�??婵犵數濮撮崐缁樻櫠濞戙垺鐓冮梺鍨儏閻忔挳鏌＄仦鍓ф创妤犵偞锕㈠鍫曞箣閻樼偣鍋℃繝鐢靛仜閻°劎鍒掑鍥ㄥ床闁告劦浜濆畷鍙夌箾閹存瑥鐏╅柣顓燁殔椤潡鎳滈悽娈跨伇闂�?€炲苯澧繛纭风�?瀵鈽夐姀鐘靛幐闂佺ǹ鏈划宥夊礆濞戞鏃堟偐闂堟稐绮跺銈嗗灥椤﹂潧顕ｉ锕€纾奸柣鎰綑閻у嫭绻濋�?锝嗙【閿燂拷?????闁哄被鍎查埛鎺楁煕鐏炲墽鎳勭紒浣哄閵囧嫰寮撮悢鍝勨拰閻庤娲忛崹浠嬪箖閸撗傛勃闁绘劦鍓氶鍥⒒娴ｅ憡璐￠柛搴涘€濋獮鎰槹鎼淬垹搴婇梺绯曞墲閵囨盯寮ㄦ禒瀣厱閻忕偛澧介。鏌ユ煕閻斿搫浠遍柡�?嬬秮楠炴﹫鎷�??閿熻棄鎲￠崚娑㈡⒑鐠団€虫灍妞ゃ劌锕顐﹀箛椤撶喎鍔呴梺鐐藉劥鐏忔瑩鎯勬惔銊︹拻濞达絿鐡旈崵娆戠磼缂佹ê鐏存鐐村姍楠炲酣鎸婃径搴㈡啺闂備胶鍋ㄩ崕杈╁椤撱垹姹查柛鈩冪⊕閸婄敻鏌ㄥ┑鍡涱€�?褌鍗抽弻銊モ槈濮橆剚鐏堝┑顔硷攻濡炰粙寮婚崨�?�樺€烽柤鑹版硾椤忣厽绻濋敓锟�?閸愩劉鎸冪紓浣介哺閹告悂顢樻總绋垮窛妞ゆ洖鎳忛敍浣虹磽閸屾瑧顦�???缂備礁顦遍幊鎾绘偩闁垮闄勭紒�?�仢�?�撳棝姊虹紒妯活梿婵炴挸�?遍懞閬嶆偨閸涘ň鎷绘繛杈剧到閹虫瑩宕烽鐔峰簥閿燂�?????闁绘挻娲熼弻娑㈩敃閿濆洤顩梺鍝勵儐閺屻劑婀�?梺缁樏Ο濠囧磿閹扮増鐓熼柟鎹愭硾閺嬫盯鏌￠敓锟�?閸犳牠寮婚崶顒佹櫇闁逞屽墴閹﹢鎮╃紒妯煎幗闂侀潧枪閸斿秹顢旈悩鐢电＜閺夊牄鍔屽ù顕€鏌熼瑙勬珔妞ゆ柨绻�?、娆撳箚瑜庨崐顖炴⒒閸屾瑧顦﹂柟纰卞亰閹绺界粙璺ㄧ崶闂佸搫绋�?崢褰掑焵椤戣法顦﹂柍璇查叄楠炴﹢寮堕幋婊勫亝闂佽楠搁崢婊堝磻閹剧粯鐓冪憸婊堝礈閻旂厧绠栭柍鈺佸暙缁剁偤鏌熼柇锕€骞愰柟閿嬫そ濮婃椽鎳￠妶鍛€炬繝銏㈡�?濡繈寮鍜佸悑濠㈣泛顑囬崢閬嶆煟鎼搭垳绁烽柛鏂跨焸閿燂拷?妞ゆ帊鑳舵晶顒傜磼�?�€鍐摵缂佺粯绻堝畷鍫曞Ω閵夈垹浜惧┑鐘崇閻撶�?鏌熼鐔风瑨闁告梹绮嶇换娑㈠川椤撶噥妫ょ紓浣介哺閹稿骞忛崨鏉戞嵍妞ゆ挻绋掗～宥嗕繆閻愵亷鎷�??閿熶粙宕�?????濞寸厧顕敓锟�????妞ゆ棁妫�??婵犳碍鐓犻柟顓熷笒閸�?鏌熷畡閭︾吋婵﹨娅ｇ划娆撳箰鎼淬垺�?�抽梻浣虹帛濡繘宕滈悢鑲╁祦闊洦绋掗弲鎼佹煥???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鎹愵嚙閻ょ偓銇勯幇鈺嬫�??閿熶粙宕瑰┑瀣厱妞ゆ劗濮撮崝婊堟煛閸涱喗鍊愰柡灞诲姂閹�?�宕掑☉姗嗕�??婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；闁绘劗鍎ら崑�?�煟濡崵�?介柍褜鍏涚欢姘嚕閹绢喖顫呴柍鈺佸暞椤忕喖姊绘担鑺ョ《闁革綇绠撻敓锟�?????缂傚倸鍊烽懗鍫曞磻閹捐纾跨€规洖娲ㄧ粈濠傗攽閻樺弶鎼愰柦鍐枑缁绘盯骞嬪▎蹇曞姶闂佽桨�?�?崯鎾蓟閵娿儮鏀介柛鈩冿供濡�?�顪冮妶蹇氱闁稿骸纾Σ鎰板箳濡や緤鎷�?閿熻姤銇勯幒鍡椾壕闂佸憡鏌ｉ崐妤冩閹炬剚鍚嬮柛婊冨暢閸氼偊鎮楀▓鍨灈妞ゎ厾鍏樺畷瑙勩偅閸愩劎鐤€婵炶揪绲介幉锟犲磹椤栫偞鈷掑ù锝呮啞閸熺偛銆掑顓ф疁鐎规洖缍婇、娑樷堪閸愩劎浜伴梻浣圭湽閸ㄥ綊骞夐敓鐘冲亗闁绘梻鍘х粻瑙勭箾閿濆骸澧�?柣蹇ｅ櫍閺屾盯鎮㈤崫銉ュ绩闂佸搫琚崝鎴�?箖閵堝纾兼繛鎴烇供閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粍顨ラ悙�?�稿ⅹ閼挎劖銇勯幒鍡椾壕婵犵鎷�??閿熷鍋㈤柡�?嬬秮楠炴帡骞嬮悩杈╅┏闂備線娼уú銈忔嫹?閿熸垝鍗抽悰顕€骞掗敓锟�??缁狅絾绻濋棃娑樻殭濞存粌澧界槐鎺炴嫹?閿熺瓔浜炲銊╂煛鐎ｎ亞效闁绘搩鍋婂畷鍫曞Ω閿旇瀚界紓鍌欒兌閿燂�??缂佺姵鐗犲璇测槈濠婂懐鏉搁梺鍝勬川閸嬫稒绂掑Ο鑽ょ瘈婵炲牆鐏濋弸娑欍亜閿曚椒鍚俊鍙夊姍楠炴帡骞樼€靛摜肖闂備線娼ф灙闁稿孩濞婇�?�鏍磼閻愮补鎷洪梻渚囧亞閸嬫盯鎳熼娑欐珷闁告挆鍛紳閻庡箍鍎遍幊蹇浰夐悙鐢电＜闁稿本姘ㄨ倴闂佸湱鎳撶€氼參骞忛崨鏉戝嵆闁绘ê寮堕悘鍫ユ⒑缁洘鏉归柛�?�尭椤啴濡堕崱妤冪懆闁诲孩鍑归崣鍐春濞戙垹绠ｉ柣妯兼暩閿涙粌顪冮妶鍡欏缂佸甯炵划鍫ュ礃椤旂晫鍘告繝銏ｆ硾閿曪妇绮斿ú顏呯厸閻忕偛澧介妴鎺楁煃瑜滈崜銊х礊閸℃稑纾婚柛娑卞灟閻掑﹥銇勯幘璺烘瀭濞存粍绮嶉妵鍕疀閹炬剚浠奸梺鍝勬４缁蹭粙鍩為幋锕€鐏崇€规洖娲ら悡鐔兼�?�鐟欏嫭�?€鐎规洦鍓濋悘鍐⒑閸涘﹤濮�?ù婊勭箞�?�曟娊顢涢悙绮规嫽婵炶揪绲块悺鏃堝吹濞嗘挻鍊垫繛鎴炲笚濞呭⿵鎷�?閿熻姤娲�?悷銊╁Φ閹版澘绠抽柟�?�稿Х閸橆剟姊绘担鍛婂暈闁告棑绠撳畷浼村冀椤愩倓绗夐梺鍝勭▉閸樹粙鎮￠妷鈺傜厽闁哄倹�?�ч幆鍫�??閿熻姤绻堥弻娑㈡倻閸℃浠稿┑顔硷攻濡炶棄鐣烽敓锟�?瀹曪絾寰勭€ｎ亜澹嶉梻鍌欒兌鏋柨鏇樺€濋垾锕€鐣￠幍顔芥闂侀潧楠忕槐鏇€€呴悜鑺ュ€甸柨婵嗛娴滄劙鏌熼柨�?�仢婵﹥妞藉畷銊︾節閸曨厾鏆ら梺璇插绾板秹骞冮崒鐐靛祦闊洦绋掗弲鎼佹�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鐗堟緲閸戠姴鈹戦悩瀹犲缂佺媭鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鍓х帛閸嬫﹢鏌曢崼婵愭Ц闁绘劕锕﹂幉姝�?�?濞戞ǹ鎽曢梺鍓插亖閸庢煡鍩涢幋鐘电＝濞达絽顫栭鍛弿濠㈣埖鍔栭悡鏇㈠箹鐎涙鈽夐柍褜鍓氱换鍫ョ嵁閸愵喗鏅搁柣妯哄暱娴滄粓姊洪崗鑲┿偞闁哄懏绋栭妵鎰板礋椤栨稈鎷洪梺纭呭亹閸嬫盯宕濋敂濮愪簻闁靛闄勫畷宀嬫嫹?閿熻姤娲樺畝鎼佸箖瑜斿畷濂稿閵忊晛鏅梻鍌欑閹测剝绗熷Δ鍛偍闁绘劦鍓氬▍蹇涙⒒閸屾瑧顦﹂柟纰卞亝瀵板嫰宕堕敓锟�?閻掑灚銇勯幒鍡椾壕缂佸墽铏庨崣鍐嚕閹惰棄骞㈡繛鎴炵懅閸樻捇鎮峰⿰鍕煉鐎规洘绮撻幃銏☆槹鎼淬垺顔曢梻浣虹帛椤ㄥ懘鎮ф繝鍥х？闁绘柨鍚嬮悡蹇撯攽閻樿尙绠抽柣锝呭船闇夐柣妯虹湴閸嬨垺鎱ㄦ繝鍛仩闁圭懓�?�版俊鎼佸Ψ閿斿彞绨存繝鐢靛У椤�?牠宕伴弽顓ф晪妞ゆ挶鍨洪崕澶嬨亜韫囨挻绁╂俊顖氬濮婃椽宕崟顓犱紘闂佸摜濮甸幐楣冨礆閹烘垟鏋庨柟鎯у暱閻庮厼顪冮妶鍡樷拹闁稿骸纾濠呫亹閹烘挴鎷绘繛杈剧到閹芥粓寮搁崘鈺€绻嗘俊鐐靛帶婵″尅鎷�?閿熻姤婢�?敃銉х紦閻ｅ瞼鐭欓悹鎭掑妿濞煎姊绘担绋款棌闁稿妫濆畷鐗堟償閵忋埄娲搁悷婊呭鐢鍩涢幒妤佺厱閻忕偟鍋撻惃鎴濐熆瑜庣粙鎾舵�?????妞ゆ劑鍨归～�?勬⒑鐎圭媭鍞虹紒顔界懇閵嗕線寮崼婵嬪敹闂佺粯鏌ㄥ璁规�??閿熻棄銈稿缁樼�??閿燂�??????閿燂�??閸曨偄鍋嶆繛瀵稿Т椤戝懘宕ヨぐ鎺撶厓鐟滄粓宕滃▎鎾崇厴闁硅揪闄勯崐鐑芥煕濞嗗浚妲撮柡�?�懇濮婃椽宕ㄦ繛鎺濅邯婵�?�爼骞栭敓锟�???娴ｅ壊娼╅柤绋跨仛濞呮粓姊虹化鏇炲⒉闁荤啙鍥ㄥ剨闁割偅绺鹃弨鑺ャ亜閿燂拷?閺嬬粯绗熷☉銏＄厱閹艰揪绲鹃弳顒勬煕閳哄绡€鐎规洏鍔戦、娆撳箚瑜嶇粭姘舵⒒閸屾瑧顦﹂柟璇х磿閹广垽宕掑┃鎯т壕婵﹩鍘介崐鎰殽閻愯尙绠婚柡浣规崌閿燂�?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧窛閿燂拷?????闁靛鍎查崳鎶芥煕椤愵偂閭柡灞剧洴椤㈡洟濡堕崨顔界槪闂備礁缍婇弨鍗烆渻閽樺娼栨繛宸簻�?�告繂鈹戦悩鎻掝仱婵℃彃鐗撳娲箰鎼淬垻鈹涚紓浣哄У閹瑰洤鐣峰ú顏勎ㄩ敓锟�???缂佸墎鍋ら弻鐔兼焽閿燂拷?楠炴﹢鏌涘▎蹇旑棦婵﹥妞藉畷顐�?礋椤掑�?�鍋愬┑鐐茬摠缁姵绂嶅⿰鍫嫹?閿熻姤绻濋崶鑸垫櫔闂�?€炲苯澧存鐐插暙铻栭柛娑卞櫘濡啫鈹戦悙鏉戠仸闁绘娲�?敓锟�????闁诡喗顨堥幉鎾礋椤掑偆妲堕梻浣告憸婵敻鎮ч悩璇参ュù锝囩《濡插牊淇婇鐐存暠妞ゎ偄绉瑰娲捶椤撶偛濡洪梺鐟版啞閹倿銆�?弮鍥ヤ汗闁圭儤鎸撮幏娲⒑閻撳寒娼熼柛濠冩礋瀵悂骞嬮悩鐢碉紲濡炪�?�姊婚崢褔顢楅姀銈嗙厸闁告稓澧楃涵楣冩懚閺嶎厽鐓曢柟鑸妽濞呭棙绻涢崼婊冨祮閿燂�??????闁绘鍋�??閸愵亞纾奸柤纰卞墮鐢爼鏌嶉挊澶樻█??闂佺粯蓱椤旀牠宕ラ崨瀛樷拻濞达綀娅ｇ敮娑㈡煕閵娾晜娑ч摶鐐寸箾閸℃ɑ鎯勯柡浣革躬閺屾盯濡烽幋婵囨拱閻庨潧鐭傚娲濞戞艾顣洪梺纭呮珪閸�?鍒掓繝姘亱闁割偅绮庣粻姘渻閵堝棗濮﹂柛瀣閻涱噣寮介鐔稿殙闂佺粯鍔曢敓锟�???闂備礁鎼ú銊︽叏闂堟稈鏋�???/pc闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺娲熼弫鍌炴偩鐏炶棄绗氶梺鑽ゅ枑缁秶鍒掗幘宕囨殾婵犲﹤鍟犲Σ鍫ユ煏韫囨洖啸闁汇倕娲娲偡閹殿喕铏庨柣搴㈠嚬閸橀箖鍩€椤掍胶鍟�???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鍓х帛閸嬨�?�鏌￠崘銊у闁稿被鍔岄埞鎴﹀磼濠婂拑鎷�?閿熶粙鏌嶈閸撱劎绮婚幘宕囨殾鐟滅増甯╅弫濠囨煏婢诡垰鍟悘鍫ユ⒑绾懏鐝柣妤冨█瀹曟椽鏁撻悩鑼槰闁荤姵浜介崝鎴澪涢悜鑺モ拻閿燂�??????濠电偞娼欏ú顓㈡晲閻愭潙绶為柟閭﹀墰閿涚喖姊洪幆褎绂嬮柛�?�噹閳诲秹鎮╃拠鑼啇闁哄鐗嗘晶浠嬪礆閻�?牄浜滈柕澶涚畳婢规﹢鏌嶇憴鍕伌鐎规洘甯掗～婵嬵敇閻愬瓨鐣奸梻鍌欒兌缁垶骞愭ィ鍐ㄧ獥闁哄稁鍘奸拑鐔兼煟閺冨伋褰掝敋闁秵鍊垫繛鎴烆伆閹达附鐓ユい鎾跺枔閿燂�??闂佸啿鐨濋崑鎾绘倶閻愬灚娅曞ù鐙€鍨崇槐鎾存媴娴犲鎽甸柣銏╁灣閸嬨�?�鐛�?幋锕€绀嬫い鏍ㄧ煯缁卞爼姊洪崨濠冨闁告瑥鍟撮幃浼村箻缂佹ǚ鎷绘繛鎾村焹閸嬫挻绻涙担鍐插幘濞差亜围闁搞儻绲芥禍鐐叏濮�?棗浜滅€规挸妫�?濞堝灝娅�?柛�?�工閿燂拷???妞ゃ垺鐟╅幊鏍煛娴ｆ劅鏇炩攽閿涘嫬浜奸柛濠冪墱閺侇喗绻濋崶顭掓�??閿熶粙鏌ㄩ弴鐑囨�??閿熺晫澹曢崸妤佺厽闁哄�?��?�ч幉鍝ョ磼閿燂拷?閸嬫挸鈹戦悩鍨毄濠殿喗鎸冲畷鎰磼濡粯鐝烽梺鍝勬川婵�?澹曟總鍛婄厽婵炲棗鑻禍楣冩⒑閹肩偛濡奸柣鏍帶椤曪絾绻濆顑┾晠鏌嶉崫鍕舵嫹?閿熻姤绂嶉悙鐑樷拺缂佸瀵у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠鐛�?幋锕€绠涢梻鍫熺⊕椤斿嫰姊绘担鍦菇闁稿﹥顨婂畷鎴﹀箻鐠囧弬锕傛煕閺囥劌鐏犵紒鐘崇洴閺屾盯顢曢敐鍡欘槰濡炪�?�楠哥粔鐟邦潖閾忓湱鐭欐繛鍡樺劤閸擃剟姊洪崫鍕櫤缂侇喗鎸绘穱濠囨偨缁嬭法顦板銈嗙墬濮樸劑顢欐繝鍥ㄢ拺闁荤喐澹嗛幗鐘电磼鐠囪尙校缂佸�?�甯楅妶锝夊礃閳圭偓瀚奸梻浣筋潐閸庡吋鎱ㄩ妶澶婃瀬闂侇剙绉甸悡鏇㈡煏婵炲灝鍔滈敓锟�?????妞ゆ梹顑欓崵娆撴煃閽樺妲搁摶锝夋⒑閸噮鍎涙繛鍏兼⒐缁绘繂鈻撻崹顔界亶濡炪們鍔岄幊姗€骞冭缁绘繈宕惰閻庮剚淇婇妶蹇曞埌闁哥噥鍨堕幃锟犳偄閼测晛褰勯梺鎼炲劘閸斿秶浜搁幍顔剧＜闁稿本鍑归崕鏃堟煛鐏炲墽鈽夐摶锝夋煕濠靛棗顏ら柟绋垮暙閿燂�?????鐎殿喖鐖煎畷婵嗏枎閹捐泛绁﹂敓锟�?????閿燂�??????闁哄洨鍋炲婵嬫煟濞戝崬鏋涢柍瑙勫灴閹晠宕归锝嗙槑濠电姵顔栭崰鏍敋椤撱垹鐒垫い鎺嶇閸ゎ剟鏌涢悩鎰佹疁???濠电偛妫欓幐濠氬煕閹达附鍋ｉ柛銉ｅ妼缁茬粯銇勯幒瀣仾闁靛洤瀚板顕€鍩€椤掑嫭鍋嬮柣妯垮皺閺嗭箓鏌熼崜浣烘憘闁轰礁顑夐弻宥堫檨闁告挻鐟╅幃楣冩倻閽樺顓洪梺缁樺姉閺佹悂鎯�?崼銉︹拺闁硅偐鍋涢崝妤呮煛閸涱喚銆掔紒顔硷躬閺佸啴鍩€椤掑嫬鐓橀柟杈剧畱閻擄繝鏌涢埄鍐炬畼濞寸姭鏅犲娲川婵犲懎顥濆銈嗗灥濞差參宕�?濡炪倖甯婇懗鍫曘€�????闁�?�屽墴楠炴牗鎷呭灞炬啺婵犵數鍋為崹鎯板綔闂佸搫顑呴柊锝夋偂椤愶箑鐐婂瀣捣钃遍梻浣哥－缁垶骞愰幖浣哥厴闁硅揪绠戦悡锟犳煕閳╁啨浠︾紒銊ょ矙濮婃椽宕妷銉愶綁鏌ｅΔ浣圭闁挎繄鍋犵粻娑㈠即閻樼绱叉繝纰樻閸ㄧ敻宕戦幇鏉跨疇婵犻潧顑嗛埛鎴︽⒑椤愩倕浠滈柤娲诲灡閺呭爼顢欐慨鎰盎濡炪倖鎸鹃崑鐐电矚閹稿簺浜滈敓锟�???缂傚秴锕濠氭偄绾拌鲸鏅╅梺闈浨归崕鏌ュ箹閹邦収娈介柣鎰典簻閻忣亜菐閸パ嶈含闁诡喗鐟╅、鏃堝礋椤撴繄妫紓鍌氬€风粈渚€顢栭崱娑樺瀭濠靛�?�鎲￠崐鍫曟煕閹伴潧鏋熼柍閿嬪灴閺屾稑鈽夊鍫濆闂佹椿鍘煎Λ婵嬪蓟閿濆绠抽柣鎰暩閺嗐倝鎮�?▓鍨灍鐟滄澘鍟撮妶顏呭閺夋垿鍞堕梺缁樻煥瀵鎷�??閿熻棄銈稿缁樻媴閸涘﹤鏆堥梺鐟版啞濡叉帡濡甸幇鏉跨闁冲搫鍠氬ú绋库攽閻樼粯娑ф繛灞傚妿缁粯銈ｉ崘鈺冨幈濠电偛妫�?ù姘瀶瑜旈弻銈夊级閹稿骸浠撮梺鍝勬湰閻╊垶宕洪敓鐘茬＜婵犲﹤瀚崹杈ㄤ繆閵堝洤啸闁稿鐩�?�鏍ㄥ緞閹邦剚鐎梺绋跨灱閸嬬儑鎷�?閿熺晫濮撮�?�璺ㄦ崉娓氼垱笑闁诲骸鐏氶悡鈥愁潖婵犳艾纾兼繛鍡樺姉閵堟澘顪冮妶鍡樼闁绘濮撮悾鐑藉閵堝棗浠奸柣蹇曞仧閸嬫挸鈻撴导�?�樷拺闁革富鍘奸崝�?�煙閹间緡妫戦柟骞垮灲瀹曞崬顪冪紒妯绘澑闂備胶枪閺堫剛鍠婂澶婄柈闁绘劗鍎ら悡鐔兼煙閹屽殶婵炲弶鎸抽弻鐔碱敊缁涘鐤�?梺杞扮劍閸旀牠骞嗛弮鍫濈伋闁肩⒈鍓欓崵顒勬⒒閸屾瑧鍔嶅┑鐐诧躬�?�劍娼忛埡鍌涙闂佺粯鍔曢悘姘讹綖閺囥垺鐓欓柣鎴炆戠亸鎵磽�?�ュ懏鍠�?柡灞炬礃缁绘盯宕归鐓庮潥闂佽崵濮村ú銊╁磻閵堝绠栨俊銈呭暞閸犲棝鏌涢弴銊ュ妞わ负鍔戦弻锝夊閳轰胶浠柣銏╁灲缁绘繈寮幇鐗堝€锋繛鏉戭儐閿燂拷?闂佽鍑界紞鍡樼閻愪警鏁囬柛蹇氬亹缁犻箖寮堕崼婵嗏挃缂佸鍓氶妵鍕敃閵忊晜鈻堥悗娈垮枛閸熷潡锝炲Δ鍛疄缂侇煉鎷�?閿熺氮h
        .fb_pause({pause_o[2],pause_o[0]}),
        .fb_interrupt(1'b0),       
//        .fb_new_pc(32'b0),
        .new_pc(new_pc_from_ctrl),

        .BPU_flush(BPU_flush),
        .pi_pc1(inst_addr1),
        .pi_pc2(inst_addr2),
        .if_pred_addr1(if_pred_addr1),
        .if_pred_addr2(if_pred_addr2),
        .inst_rreq_to_icache(inst_rreq),
        .pi_is_exception(pi_is_exception),
        .pi_exception_cause(pi_exception_cause),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹寸偛顥氶柛娆忔惈閳规垿鎮╅崹顐ｆ瘎婵犳鍠氶崗姗€濡撮崒娑氼浄閻庯綆浜為ˇ顓炩攽閻樼粯娑фい鎴濇噽缁寮介鐔哄幈闁诲繒鍋涙晶浠嬪煟閵壯呯＜閻犲洤寮堕ˉ銏ゆ煛瀹€瀣М妤犵偛顑夐弫鎰板川閸涱喗宕岄柡宀嬬節瀹曘劑顢欓崜褏鍘掔紓鍌欐祰妞存悂骞愭繝姘闁告稑鐡ㄩ崕�?€绱掔€ｎ亞浠㈢憸鏉挎閳规垶骞婇柛濠冾殕閹鳖煉鎷�?閿熻棄鎲″畷鍙変繆椤栨瑨顒熸繛鍏肩墱缁辨挻鎷呴懖鈩冨灦閸掑⿵鎷�?閿熻棄鎽滅壕鍏肩箾閹寸儑渚涢柛搴＄箲缁绘盯宕奸銏犵缂備浇椴搁幐濠氬箯閸涘瓨鎯為柣鐔稿椤愬ジ姊绘担鍛婂暈婵﹤缍婇妴鍐╃�?閸モ晛绁﹂梺纭呮彧缁犳垿锝為崨�?�樼厪闁割偅绻冮崵鍥煕閻愯尙鍩ｆ慨濠冩そ濡啫鈽夋潏銊愩�?�姊虹粙鍨劉濠电偛锕ㄥΛ鐔奉渻閵堝棙纾甸柛�?�尰閹便劍绻濋崨顕呬哗濠电偞鍨归弫璇茬暦閵娾晩鏁婇柛蹇撱偢閺侇亝绻濋悽闈浶ユい锝勭矙閿燂拷?妞ゆ帒鍟悵顏堟煙閸忕厧濮嶉柡宀嬬秮閺佹劙宕堕妸锔界槗闂備浇妗ㄩ悞锕傚箲閸ヮ剙鏋�?柟鍓х帛閺呮悂鏌�???闂傚倸鍊烽懗鍓佸垝椤栫偛绠归柍鍝勬噹绾捐鈹戦悩璇ф嫹?閿熶粙寮抽敃鍌涚厱妞ゆ劧绲鹃敓锟�??闁诡垳鍠栭幃宄扳堪閸愮偓效闂�?€涚┒閸�?垵鐣烽崼鏇ㄦ晢濞达絽寮剁€氳偐绱撻崒娆戭槮妞ゆ垵妫濋、鏍р枎閹惧磭锛熷┑鐐村灦閳笺倝鎮�???闂佸憡娲﹂崢楣冩偪閸曨剛绡€缁炬澘顦辩壕鍧楁煛娴ｇ瓔鍤欓柣锝囧厴閹垻鍠婃潏銊︽珫婵犳鍠楅敃鈺呭礈濞嗘挸鏋�?柕鍫濐槹閳锋帒霉閿濆懏璐￠敓锟�?娴犲鐓曢柕濞垮妽椤ュ銇勯鐐寸┛閿燂�??????闁哄洠鍓濋鐘裁归悪鍛洭闁瑰弶鎸抽弫鎰板幢濡粯绶梻鍌氬€烽懗鍓佸垝椤栫偛绀夋俊顖炴？閻掑﹥绻涢崱妯哄婵炲懐濞€濮婃椽顢�?缂佸鏁婚幃锟犲即閵忥紕鍘繝鐢靛仜閻忔繃淇婇悾�?€妫い鎾跺Т娴滈箖鏌曢崶褍顏い銏℃礋閿燂拷?闁靛繈鍩勯崬铏圭磽閸屾瑦绁板鏉戞憸閺侇噣骞掗弴鐘辫埅闂備浇宕垫慨鏉懨洪妶鍛傜喐绻濋崶褏鍔﹀銈嗗笂閻掞箑鐣风仦鐐弿濠电姴鍟妵婵撴嫹?閿熻姤娲�?〃濠傤潖閼姐倕顥氶悗锝庝簽閸旂敻姊婚崒娆掑厡?闁诲孩绋堥弲婊呮崲濞戞瑧绡€闁告剬鍛暰闂佽�?�╃粙鎺椻€﹂崶鈺佸К闁�?�屽墴濮婃椽骞栭悙鎻掑闂佸憡鏌ㄩˇ鐢哥嵁韫囨拋娲敂閸涱亝�?�奸梻浣告啞缁嬫垿鏁冮敂鍓х＝婵ǹ鍩栭悡鏇㈠箹濞ｎ剨鎷�??閿熶粙宕ú顏呯厽??闂佸府绲介～蹇曠磼濡顎撻梺鍛婄☉閿曘倝寮抽崼婵冩�?妞ゆ梻銆嬪銉х磽瀹ュ拑韬鐐插暣閹粓鎸婃竟鈹垮姂閺屽秹宕崟鑸垫暰闂佸搫鎷嬫禍顏勵潖濞差亜绠伴幖杈剧悼閻ｉ潧顪冮妶蹇撶槣闁搞劋鍗抽�?�娆掔疀閹绢垱鏂€闂�?潻鎷�??閿熺晫绠�???闂傚倷鑳剁划顖濇懌閻熸粍婢橀崯鎾€�?弮鍫晝闁挎梻鏅崢浠嬫⒑閹稿孩纾甸柛�?�崌閿燂拷???婵☆偅绻堝畷娲倷閸濆嫮顓洪梺鎸庢⒒缁垶寮查埡鍛拺閿燂拷?????闂佺ǹ锕ラ幐鎯р枎閵忋�?�鍋ㄩ柛娑樑堥幏娲⒑閸涘﹦鈽夐柨鏇樺劤娴滃憡�?�肩€涙鍘介梺鍐叉惈閿曘�?�鎮�?敃鍌涚厪闁糕剝娲滈ˇ锕傛煃鐠囨煡鍙勬鐐达耿�?�曟﹢鎳犻崹娑樹壕闁割煈鍠掗弨浠嬫煟閹邦厽缍戦柣蹇ョ畵閺岋綁鎮㈤弶鎴犱紙濡ょ姷鍋涚换妯虹暦椤愶箑�?嬮敓锟�????濠碉紕鍋戦崐鏍ь潖婵犳艾纾婚柟鎹愵嚙閸氬綊鏌嶈閸撴瑩鍩為幋锔藉€烽柤纰卞墯閸曢箖姊虹粙鍖℃敾缂佽鐗嗛悾宄懊洪鍕姦濡炪�?�甯婇梽宥嗙濠婂牊鐓欓悗鐢登规禒锕傛�?�濮橆厽�?嬮柡�?€鍠栧畷娆撳Χ閸℃浼�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牗绋戞禒濂告⒑濮瑰浄鎷�??閿熶粙宕归浣侯洸鐟滅増甯楅悡娆撴煟閹寸倖鎴犱焊閻㈠憡鐓曢柡鍌濇硶閸╋綁鏌熼绛嬫畼闁瑰弶鎸抽敓锟�???闁藉嫬銈稿铏圭矙閸ф寮版繛瀛樼矋閸庣厧螞閻斿娓婚柕鍫濇婢ч亶鏌涚€ｎ偆娲撮柟顕嗘�??閿熻В�?介悗锝庝簽椤�?劕鈹戦悜鍥╃У闁告挻鐟︽穱濠囨嚃閳哄啰锛滈梺缁樏幖顐�?触閸︻厾纾奸弶鍫涘妼濞搭喗銇勯姀锛勬噧闁宠閰ｉ幃娆擃敆閸屾簽銉╂⒒娴ｇ瓔鍤欓悗娑掓櫊閹虫繃銈ｉ崘銊幯呯磼鐎ｎ偒鍎ユ繛鍏肩墬缁绘稑顔忛鑽ゅ嚬闂佹悶鍊栫敮锟犲蓟閺囥垹閱囨繝闈涙搐閺呬粙姊洪幐搴ｇ畵闁诡喖娼￠幃鐑藉箥閸愯尙澧梻渚婃嫹?閿熻棄鑻晶浼存煕閹烘挸绗掗柍璇叉唉缁犳盯寮撮悢鍓插晭濠电姷鏁搁敓锟�??婵炰匠鍥ㄥ亱闁告侗鍘搁弻锔姐亜韫囨挾澧涢柛�?�у墲缁绘盯宕卞Ο鍏煎櫘缂備礁顑呴�?�鐑藉蓟閿濆棙鍎熼柕寰涢铏庢繝娈垮枛閿曘劌鈻嶉敐澶婄疅闁圭虎鍠栫粈瀣亜閹伴潧浜濇い銉ヮ儏閳规垿鎮╅锝咁€忛梺鍛婃礀閻忔岸鎮块敓锟�?閹鈻撻崹顔界亶闂佺粯鎼换婵嬫偘閿燂�??瀵粙濡搁敓锟�?椤庢捇姊洪棃鈺佺槣闁告鍘ч锝夊箮閼恒儮鎷绘繛杈剧秬濞咃絿鏁☉娆戠闁告瑥顦辨晶纰夋嫹?閿熻姤娲�?崝姗€濡甸幇鏉跨闁规儳鐡ㄩ鐔兼⒒娴ｈ姤纭堕柛锝忕畵閿燂拷??????
        .ex_is_bj(ex_is_bj),
        .ex_pc1(ex_pc1),
        .ex_pc2(ex_pc2),
        .ex_valid(ex_valid),
        .real_taken(ex_real_taken),
        .real_addr1(ex_real_addr1),
        .real_addr2(ex_real_addr2),
        .pred_addr1(ex_pred_addr1),
        .pred_addr2(ex_pred_addr2),
        .get_data_req(get_data_req),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹瑩寮堕崹顕呭殭闂傚�?�鍊搁崐鐑芥倿閿曞�?�绠栭柛顐ｆ�?绾惧潡鏌ｉ幋鐑嗙劷妞も晛寮剁换婵囩節閸屾粌顤€闂佺ǹ楠哥粔褰掑蓟閿濆绠ｉ柣鎰�?暞缁秶绮嬪鍛牚闁割偆鍠撻崣鍡涙⒑閸濆嫬鏆欐繛鏉戝€垮畷闈涒枎閹存柨浜炬繛鍫濈仢濞呮﹢鏌涢敐蹇曠М鐎殿喖顭烽崹鎯х暦閸ャ劍鐣烽梺璇插嚱缂嶅棝宕滃☉婧惧徍闂傚倸鍊峰ù鍥敋閺嶎厼绐楅柟鐑橆殔閻ょ偓绻濇繝鍌氭灓闁绘帊绮欓悡顐﹀炊閵娿�?�绻�?梺杞扮閸燁垶濡甸崟顖氱�?闁宠桨鑳舵禒濂告⒒婵犲繒鐣垫慨濠傤煼瀹曟帒顫濋钘変壕闁绘垼濮ら崵鍕煕閹捐尙顦﹂柛銊︾箖閵囧嫰寮介顫捕缂備胶濮抽崡鎶藉蓟閻斿吋鈷掗悗鐢登规俊浠嬫⒑缁嬫鍎忔い鎴濐�?瀵鎮㈤崗纭锋�??閿熻姤銇勯幒鍡椾壕婵犫拃灞界仸闁哄本鐩俊鍫曞幢濡⒈妲归梻浣告惈閺堫剟鎯勯鐐靛祦闁搞儺鍓﹂弫鍥煟濮�?棗鏋涘ù鐙呯畵濮婄粯鎷呯粙娆炬闂佺ǹ顑嗙敮妤冪矉�?�ュ鏁傞柛顐ｇ箚閹芥洖鈹戦悙鏉戠仧闁糕晛�?�板顐�?礃椤旂晫鍘梺鍓插亝缁诲啴宕冲ú顏呯厽闊洤娴风粣鏃€鎱ㄦ繝鍐┿仢鐎规洏鍔嶇换娑㈠箳濠靛懘鍋楅梺璇″枟閿氭い顐ｇ箞椤㈡﹢鎮╅锝嗘殼婵犵數濮烽弫鍛婃叏閺夋嚚娲晝閸屾氨锛欐俊鐐差儏缁ㄥ爼宕戦幘缁樺仭闁哄顑欏Λ宀勬⒑閸濄儱校闁绘濮撮悾宄扳堪閸喎浜遍梺鍓插亝缁海绮诲鑸碘拺闂傚牊绋撴晶鏇熺箾鐏炲偊鎷�??閿熶粙鎮ф惔銊︹拻濞达絿鐡旈崵鍐煕閻樺磭澧电€规洘鍔欓獮鏍ㄦ媴閻熼鎮ｉ梻浣虹帛閸ㄧ厧螞閸曨垽缍栭柛娑樼摠閻撳繘鏌涢锝囩畺闁革�?濮ら敓锟�????閻㈩垱甯￠垾鏃堝礃椤斿槈褔鏌涢埄鍏︽岸骞忔繝姘拺闁告繂瀚刊濂告煕鐎ｎ亷宸ラ柣锝囧厴閿燂拷?闁靛牆鎳庣粣娑欑�?閻㈤潧孝閻庢凹鍣ｉ�?�娆撳即閵忥紕鍘告繝銏ｆ硾閿曪附鏅堕弴鐑嗙唵鐟滃繘寮查銈呭灊闁哄啫鐗滈弫鍡椕归敐鍛�?�缂併劏顕ч�?�鍐Χ閸℃顫囬梺绯曟櫅鐎氼剙宓勯梺褰掓？閻掞箓鎮￠悢鍏肩叆婵犻潧妫欓崳瑙勪繆閹绘帩鐓奸柡宀嬬秮閺佹劙宕卞▎鎴犳澖闁诲氦顫夊ú婊堝窗閺嶎叏鎷�?閿熻棄螖閸涱厾锛滃┑顔斤供閸撴盯顢樻總鍛娾拻閿燂�??????闂佺粯甯粻鎾崇暦閺囥垹�?冮悷浣疯兌閹虫捇锝炲┑鍫熷磯闁惧繒娅㈢槐顕€姊虹拠鎻掑毐缂傚秴妫濆畷鎶筋�??鐎殿噮鍋婂畷鎺楁倷鐎电ǹ骞堟俊鐐€栭崝锕傚磻閸曨剚娅犻柟娈垮枤绾惧ジ鎮楅敐搴濈敖缂佺姳鍗抽弻宥囨喆閸曨偆浼岄梺璇″枓閺呮繄妲愰幒鎳崇喐绻濆顓熸婵犵绱曢崑鎴�?磹閺嶎厼鍨傞柣銏⑶圭粻鐘绘煙闁箑鍘存俊鎻掔墦閺岋綁濮€??闂佺粯甯掗悘姘跺Φ閸曨垰绠抽柟瀛樼箥娴犻箖姊洪幎鑺ユ暠闁搞劌婀卞Σ鎰板箻鐎涙ê顎撴繝娈垮枟閸╁牊绂嶅┑瀣疄闁靛ň鏅涢悙濠冦亜閹哄秷鍏岄柛妯圭矙濡懘顢曢姀鈥愁槱闂佸搫琚崝鎴濈暦椤愶附鍊绘俊顖炴櫜缁ㄥ姊洪棃娑氱畾闁糕晛�?�伴獮�?�偐閸愭彃绨ユ繝鐢靛█濞佳兾涢鐑嗙劷闁冲搫鍊舵禍婊堟煙閹屽�??闂佽�?�╂穱鍝勎涢崟顖氱厴闁硅揪闄勯崐鐑芥煠閹间焦娑ф繛鎳峰懐纾藉ù锝囨嚀缁茬粯绻�?????闁伙絿鍏樺鎾閻樻爠鍐剧唵閻犺櫣灏ㄥ銉╂煙椤栨粌浠辨慨濠冩そ閺屽懘鎮欓懠璺侯伃婵犫拃鍐憼闁�?�究鍔嶇换婵嬪礃閳瑰じ铏庢俊銈囧Х閸嬬偤鎮ч悩璇茬畺婵犲﹤鐗嗛悙濠囨煏婵炲灝鍔撮敓锟�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楃€广儱娲ら崹婵囩箾閸℃ɑ灏紒鐘崇墱閹叉悂寮崼婵堢暫闂佸啿鎼崯顖ゆ�??閿熻姤宀搁弻娑樷枎韫囷絾楔闂�?€炲苯澧婚柛鎾跺枎椤繐煤椤忓懎浠梺鍝勵槸缁ㄩ亶骞愰崘顏嗙＝濞撴艾娲ゅ▍姗€鏌涢妸銊︾【妞ゆ洩缍佸濠氬Ψ閵壯屽晣濠电偠鎻徊钘夛�?�闁�?秴鐭楅柛鈩冪⊕閳锋垹绱撴担鐧告嫹???闂備胶枪閿曘倕锕㈤柆宥呯劦妞ゆ帊鑳堕崯鏌ユ煙???
        .fb_pred_taken1(fb_pred_taken1),
        .fb_pred_taken2(fb_pred_taken2),
        .fb_pc_out1(fb_pc1),
        .fb_pc_out2(fb_pc2),
        .fb_inst_out1(fb_inst1),
        .fb_inst_out2(fb_inst2),
        .fb_valid(fb_valid),
        .fb_pre_branch_addr1(fb_pre_branch_addr1),
        .fb_pre_branch_addr2(fb_pre_branch_addr2),
        .fb_is_exception1(fb_is_exception1),
        .fb_is_exception2(fb_is_exception2),
        .fb_pc_exception_cause1(fb_pc_exception_cause1),
        .fb_pc_exception_cause2(fb_pc_exception_cause2),
        .fb_instbuffer_exception_cause1(fb_instbuffer_exception_cause1),
        .fb_instbuffer_exception_cause2(fb_instbuffer_exception_cause2)
    );


    backend u_backend(
        .clk(aclk),
        .rst(rst),

        // from outer
        .is_hwi(intrpt),
        
        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儵姊婚崒娆掑�??闂佹寧娲忛崐婵嬪灳閿燂拷?閻ｏ繝鏌囬敓锟�?濞堛劑姊虹憴鍕姸濠殿喓鍊濆鎻掆堪閸喓鍘介梺鎸庣箓閹虫劙鎮橀柆宥嗙厽??闁绘锕﹂幑銏犫攽鐎ｎ偄浠洪梻鍌氱墛閿燂�??闁靛繈鍊栭悡鏇炩攽閻樻彃鏆為敓锟�??????妞ゆ棁濮ら崐鎰攽闄囬崺鏍ь嚗閿燂�???閿濆骸澧鐐茬墛缁绘繂鈻撻崹顔界亶闂佹寧娲嶉弲鐘茬暦濠婂牊鏅濋柛灞炬皑閿涚喖妫呴銏�?�闁哄矉绲剧粋宥呪堪閸曗晙绨婚梺鍦檸閸ㄧ増鏅堕懠顒傛／妞ゆ挾鍋熼崺锝夋煛閿燂�??閸犳牠骞冮悜钘夌骇婵炲棗褰為�?顏嗙磽閸屾瑧鍔嶆い銊ョ墦瀹曚即寮�?????濠电偞鍨堕敃鈺侇焽閳哄�?�浜滈柟鍝勬娴滄儳顪冮妶鍐ㄥ姎濡ょ姵鎮傞崺鐐哄箣閿旇棄浜归梺鍓茬厛閸嬪懎袙閸曨垱鈷戠紒瀣儥閸庢劙鏌ｉ埡濠傜仸闁绘侗鍠楃换婵嬪磼濠婂嫭鐣烽梻浣告啞濞诧箓宕戦崟顖涘€垫い鎾卞灪閳锋垿鏌ら幁鎺戝壄妞ゅ繐鐓婚崶顒佸癄濠㈣埖顭囬崝鐑芥⒑閸濆嫮袪闁告柨娴风划濠氬礈瑜夐崑鎾绘偡閺夋妫岄梺鍝ュУ濞叉粓鎳為柆宥嗗殥闁靛牆鍊告禍楣冩煟閻斿搫顣奸柛鐔哄仧缁辨帞鎷犻敓锟�???閸ф鏄ラ柣鎰惈缁狅綁鏌ㄩ弮鍥棄濞存粌缍婂娲捶椤撶姴绗￠柣銏╁灡椤ㄥ懘鍩㈤幘娲绘晣闁绘鏁搁敍婊勪繆閵堝繒鍒伴柛鐕佸灦瀵啿饪伴崼鐔哄幐闂佸憡渚楅崰姘洪幘顔界厱闁冲搫鍟禒杈殽閻愬樊鍎旈柡浣稿€块幐濠冨緞閸℃ぞ澹曟俊鐐差儏缁ㄥ爼宕戦幘缁樺仭闁哄顑欏Λ�?勬⒑閸濄儱校妞ゃ劌妫濆鏌ュΨ閵夈垺鏂€闂佺粯锚閻忔岸寮抽埡鍛厱閻庯綆鍓欏暩婵炲瓨绮庢灙闁宠閰ｉ獮妯虹暦閸モ晛鐐婇梻鍌欑閹碱偆绮旈弻銉ョ閻庯綆鍓氬畷鏌ユ煕閳╁啰鈯曢柣鎾寸懅缁辨挻鎷呴棃娑氫患闂佸搫顑嗙粙鎾绘儉椤忓牆绠氱憸�?�磻閵忋�?�鐓涢敓锟�?鐎ｎ剛袦濡ょ姷鍋涘ú顓€€佸Δ鍛＜婵炴垶鐟ラ弸娑樷攽閻樺灚鏆╅柛�?�洴楠炲﹤鐣濋崟顐㈢€梺鑺ッˇ钘夘焽閺嶎厽鐓ｉ煫鍥ㄥ嚬濞兼劧鎷�?閿熻姤娲栭ˇ鐢稿蓟閺囩喓绠鹃柛顭戝枛婵洟姊虹紒妯肩細闁搞劏妫勯～蹇撁洪鍛画闂佸搫顦伴敓锟�????闂傚倷鑳堕幊鎾诲吹閺嶎厼绠�???婵犵數濮烽弫鍛婃叏閹绢喗鍎夊鑸靛姇缁狙囧箹鐎涙ɑ灏ù婊呭亾娣囧﹪濡堕崟顓炲闂佸憡鐟ョ换姗€寮婚敐澶婄闁挎繂妫Λ鍕磼閹冣挃缂侇噮鍨抽幑銏犫槈閵忕姷顓洪梺缁樺姈椤旀牠寮抽敓鐘冲€甸悷娆忓閿燂�??閻庢鍠栭悥濂哥嵁閸儱惟闁靛鍠楃€靛矂鏌ｉ悩鍙夌┛鐎殿喗鎸荤粩鐔煎即閻斿墎绠氶梺闈涚墕濞层�?�鏆╅梻浣呵归鍡涙儎椤栨氨鏆︽い鏍剱閺佸啴鏌ㄩ弬鎸庢儓濞存粌鍚嬬换娑㈠级閹存繃鍊┑鐐插悑閻熲晠寮荤€ｎ喖鐐婃い鎺嶈兌閸樹粙姊洪崫鍕殭闁绘锕顐︽焼�?�ュ棛鍘介梺闈涚墕閹冲繘宕甸崶銊�?弿濠电姴瀚敮娑氱磼濡ゅ啫鏋�???濡炪倖宸婚崑鎾淬亜椤撶偞绌挎い锕€缍婇弻鈩冩媴鐟欏嫬纾抽梺杞扮劍閹瑰洭寮幘缁樻�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柛婵勫劗閸嬫挸顫濋悡搴☆潾闂�?€炲苯澧柣顓у櫍瀹曪繝骞庨挊澹┿儱銆掑锝呬壕閻庢鍣崳锝呯暦婵傚憡鍋勯柧姘€婚惄搴ㄦ⒒閸屾瑨鍏�??缂備胶绮崝娆撳箚閸愵喗鍊婚柦妯侯槺椤斿棛绱撻崒娆戝妽妞ゎ厼娲ㄧ划缁樸偅閸愩劎楠囬梺鍓插亝缁诲�?�鍩涢弮鍫熺厱闁瑰搫绉村畵鍡涙煛閿燂�??閸犳捇宕版繝鍥х闁绘劖澹嗛弫鏍⒒娴ｈ姤銆冪紒璁圭節瀹曟娊鏁愰崨顖涙婵犻潧鍊绘灙闁告濞婇弻锝夊棘閹稿孩鍎撳Δ鐘靛仦椤ㄥ﹤顫忓ú顏勬嵍妞ゆ挾鍋涙俊鐑樼�?閻㈤潧浠滈柨鏇樺€濋幃鎯х暋閹佃櫕鏂€闂佺硶鍓濋悷锕€鈻撻弴銏�?拺闁告稑锕ラ敓锟�??婵犫拃鍐╂崳缂侇喗鐟ㄧ粻娑㈠箻椤栨稒鏉搁梻浣虹帛椤洨鍒掗姘ｆ鐟滃酣濡甸崟顖氱婵犻潧娲ゅ▍銈夋⒑缁嬪灝鐦ㄩ柛�?�躬�?�鏁愭径瀣簻闂佸憡绺块敓锟�????闂傚倷鐒�?鍧�?储婵傜ǹ纾归柛褎顨堝畵渚€鏌涢幇闈涙灍闁稿﹦鍏�?幃妤呮濞戞瑦鍠愰梺浼欑畱閻楁挸顫忓ú顏勭闁绘劖褰冩慨宀勬⒑閸涘﹥鐓ラ梺甯到閻ｇ兘濮€閵堝孩鏅滈梺鍛婁緱閸ㄦ娊鎯侀崼銉︹拺婵懓娲ら悘鍙夌箾娴ｅ啿瀚々椋庢喐閺冨牆钃熸繛鎴炲焹閸嬫捇鏁愭惔鈥茬凹闁诲繐娴氶崣鍐蓟�?�ュ洦�?�氶柤纰卞劮????闁哄洦锚婵倹銇勯姀锛勨�??闂佸憡绮岄崯鐗堟償婵犲洦鈷掗柛灞剧懆閸忓瞼绱掗鍛仸闁诡喚鍏橀敓锟�??闁靛牆鎳愰敍娑㈡⒑閻熸澘鈷旂紒顕呭灦閹繝寮撮姀锛勫帾婵犵數鍋涢悘婵嬪礉閵堝鐓曢柍鍝勵儑閹ジ鏌嶈閸撴岸顢欓弽顓為棷??鐎规洘鍨剁换婵嬪炊閳轰胶銈︽繝纰樻閸ㄧ敻宕戦幇顔碱棜闁稿繘妫跨换鍡樸亜閺嶃劎鐭岄悽顖涚⊕閵囧嫯绠涢弴鐐寸亪濠殿喖锕︾划顖炲箯閸涘瓨鍤嶉敓锟�??????闂傚倷绶氬鑽ょ礊閸モ晝涓嶉柟鎹愵嚙閺嬩線鏌熼崜褏甯涢柡鍛倐閺屻劑鎮�??????
        .new_pc(new_pc_from_ctrl),
        .pc_i1(fb_pc1),
        .pc_i2(fb_pc2),
        .inst_i1(fb_inst1),
        .inst_i2(fb_inst2),
        .valid_i(fb_valid),
        .pre_is_branch_taken_i({fb_pred_taken2,fb_pred_taken1}),
        .pre_branch_addr_i1(fb_pre_branch_addr1),
        .pre_branch_addr_i2(fb_pre_branch_addr2),
        .is_exception1_i(fb_is_exception1),
        .is_exception2_i(fb_is_exception2),
        .pc_exception_cause1_i(fb_pc_exception_cause1),
        .pc_exception_cause2_i(fb_pc_exception_cause2),
        .instbuffer_exception_cause1_i(fb_instbuffer_exception_cause1),
        .instbuffer_exception_cause2_i(fb_instbuffer_exception_cause2),

        .bpu_flush(BPU_flush),   // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佸憡鏌ㄧ粔璺衡槈閻㈠憡鍊锋い鎴濆綖缁ㄨ顪冮妶鍡楀闁搞劏宕电划缁樺鐎涙ê浜楅梺闈涚墕濡孩绂嶅⿰鍫㈠彄闁搞儯鍔嶇亸顓熴亜韫囧﹥娅婇柡�?嬬稻閹棃顢欓悡搴ｎ啇婵＄偑鍊ゆ禍婊堝疮鐎涙ü绻嗛柛顐ｆ礀楠炪垺淇婇婧炬嫛婵″樊鍓熷缁樻媴閻戞ê娈岄梺鍝ュ枎濞硷繝寮绘繝鍥ㄦ櫜闁告侗鍨卞▓鎯р攽閻樿宸ラ柣妤€锕幃鐐烘嚃閳规儳浜炬鐐茬仢閸旀碍淇婇銏㈢劯妤犵偛绻愮叅妞ゅ繐鎳夐幏娲⒑閸涘﹦鈽夐柨鏇缁骞樼紒姗堟嫹?閿熻姤鎱ㄥΟ鐓庡付鐎殿噮鍣ｉ幐濠囨偄閸忚偐鍘介梺褰掑亰閸犳寮抽埡鍐／闁诡垎鍐╁€梺闈涙搐鐎氭澘顕ｉ敓锟�?瀹曟儼顦辨慨瑙勵殜濮婅櫣绱掑Ο铏诡儌閿燂拷????鐎殿喖顭烽弫鎰板醇閵忋垺婢戦梻浣烘嚀閻忔繈宕锕€�?堥悹楦裤€€閺€鑺ャ亜閺冨偊鎷�?閿熶粙寮ㄧ紒妯圭箚闁绘劘鍩栭ˉ澶愭煟閿濆洤鍘存い銏℃礋閺佸啴鍩€椤掑�?�鐭嗛悗锝庡枟閻撴洘銇勯鐔风仴闁�?�屽墾缂嶄線寮崘顔肩＜婵炴垶甯楃€氬ジ姊洪懡銈呅㈡繛娴嬫櫇娴滅ǹ鈻庨幋鐘辩瑝闂佽偐鈷堥崜娑氬婵傚憡鍋ｉ柛銉簻閻ㄥ搫顭胯缁犳捇寮婚弴銏犲耿闁哄洨濮烽悰銏ゆ�?�濞堝灝娅橀柛锝忕到閻ｉ攱绺介崜鍙夋櫇闂佹寧绻傚Λ娆撴偟濠靛鈷掗柛灞剧懅缁愭梹绻涙担鍐插濞堜粙鐓崶銊︾妞ゎ偅娲熼弻锟犲炊閵夈儳浠奸梺绋胯閸旀垿寮诲☉妯锋婵鐗嗘慨娑氱磽娴ｅ搫鈻堢紒鐘崇墪椤曪綁宕奸弴鐐哄敹濠电�?娼уΛ宀勫箰閸愵亞纾藉ù锝呭濡牓鏌涢幘鏉戝摵濠碉紕鏁诲畷鐔碱敍閿濆棙娅囬梻渚€娼х换鍡涘疾濠婂懐鎳呴梻鍌氬€峰鎺旀椤�?儳绶ゅù鐘差儏鎼村﹪鏌＄仦璇插姕闁稿鏅滅换婵嬫濞戝崬鍓伴梺缁樺笒閻忔岸濡甸崟顖氱闁瑰瓨绻嶆禒濂告⒑缂佹ê绗掗柣蹇斿哺婵＄敻宕熼姘鳖唺閻庡箍鍎卞ú鈺冪玻濡ゅ懏鈷戦柛婵勫劚閺嬪海绱掔紒姗堣€跨€殿喛顕ч埥澶愬閳╁啯鐝抽梺纭呭亹鐞涖儵宕滃┑瀣仧婵犻潧顑嗛崐鐢告偡濞嗗繐顏敓锟�?閸愵亞纾兼い鏃囧Г瀹曞本顨ラ悙鎻掓�???闂侀潧鐗嗗Λ宀勫箯瑜版帗鈷戠憸鐗堝笒娴�?即鏌涢悩鍐插摵闁诡喚鍋撻妶锝夊礃閳圭偓�?�藉┑鐐舵彧閿燂�???濡炪們鍎辩换姗€寮�????妞ゅ繐鎳庡▍锝夋煟閹炬唻鎷�?閿熶粙寮婚垾鎰佸悑閹艰揪鎷�?閿熺晫顔�????闁规崘灏欑粣鏃堟煛鐏炵偓�?夌紒鐘崇⊕缁绘盯骞嗚婢规洟姊洪懖鈹炬嫛闁告挻鐩幃鐐偅閸愨斁鎷绘繛鎾村焹閸嬫挻绻涙担鍐叉处閸嬪鏌涢埄鍐槈缂佺媭鍨堕弻鐕傛�??閿熻姤顭囩粻銉︾箾閸忚偐澧ǎ鍥э躬婵�?�爼宕ㄩ鐔割啀缂備胶鍋撻崕鎶藉Χ閹间礁钃熼柣鏃傚帶缁犵敻鏌熼悜妯肩畵闁告挻濞婂鐑樺濞嗘垵鍩岄梺璇茬箲瀹€鎼佺嵁閸儱惟閿燂拷????闂備胶枪鐞氼偊宕愬Δ鍛Е閻庯綆鍠楅崐鐢告偡濞嗗繐顏敓锟�?閸愵喗鍋ㄦい鏍ㄧ☉濞搭噣鏌涢埞鍨仾闁诡垱妫冩俊鎼佸Ψ瑜忛弶鍛婁繆閻愵亷鎷�??閿熶粙寮婚妸鈺佺妞ゆ劧绲块々鐑芥煙閻戞ê鐏嶉敓锟�??娴犲鐓熸俊顖濇娴犳盯鏌￠崱蹇�?珚閿燂拷?????妞ゆ劑鍊栭崚娑㈡煢濡崵绠為柡灞稿墲瀵板嫸鎷�??閿熻棄澧庣粚鍨攽閻愬弶鈻曞ù婊勭箞�?�曟垿宕熼顐ｅ�????妞ゅ繐�?�烽崝澶娾攽閻愯尙澧㈤柛瀣尵閹广垹鈽夐�?鐘甸獓闂佺懓鐡ㄩ敓锟�?????濠电姷鏁搁崑娑㈠触鐎ｎ喗鍋＄憸蹇涘礆閹烘梹�?�氭繛鏉戭儐椤秹姊洪棃娑㈢崪缂佽鲸娲熷畷銏ゅ川婵犲嫮鐦堥梺闈涢獜缁插墽娑垫ィ鍐╃叆闁哄浂浜顔剧磼閸屾稑娴敓锟�???闂侀潧鐗嗗Λ娑㈠储闁秵鈷戦梻鍫熺〒婢ф洘淇婇锝庢疁闁诡喗锕㈤弫鍌炲礈瑜忛敍婊呯磽閸屾瑧鍔嶆い顓炴川缁鎮欓悜妯煎幍濡炪倖妫佸畷鐢告儗濞嗘劒绻嗘い鎰╁灩閺嗘瑩妫佹径鎰仯濞达絽鎲＄拹锛勭磼婢舵ê娅嶉柡宀嬬磿娴狅妇鎷犲ù�?�壕婵犻潧顑呯粻鏍煟閹达絾顥夌紒鐙欏洤绠归悗娑櫳戠亸浼存倵閸偆澧辩紒杈ㄦ崌瀹曟帒鈻庨幋锝囩崶闂備礁鎽滄慨鐢告偋閻樿鐏抽柨鏇炲€归崐璇测攽椤旇棄濮€闁稿鎸婚幏鍛寲閺囩噥娼旈梻渚€娼х换鍡涘焵椤掍焦鐏遍柛�?�崌閹粓鎳�????闂備焦鐪归崹璇测枍閵夈劊浜归柟鐑樻煥缁侊箑鈹戞幊閸婃洟骞婅箛娑樼厱闁圭儤鍤氳ぐ鎺撴櫜闁告洦鍣�?崝鍛存⒑鐞涒€充壕婵炲鍘ч悺銊╂偂濞嗘劗绠鹃柤濂割杺閸炶櫣绱掗妸褎娅曢柍褜鍓欓悘姘熆閿燂拷?閺佸啴顢旈崟顓熸闂佽澹嗘晶妤呭磻閸℃褰掓晲閸偅缍堥梺浼欒缂嶄礁顫忔繝姘＜婵﹩鍏�?崑鎾诲箹娴ｅ摜锛欐俊鐐差儏濞寸兘鎯岄崱妤嬫嫹?閿熻棄顫濋敐鍛婵°倗濮烽崑鐐烘偋閻樹紮鎷�?閿熶粙寮撮姀鈩冩珖闂�?€炲苯澧扮紒顔碱煼閹晠鎳￠妶鍛导闂備焦鎮堕崕顖炲礉鎼淬劌鐓�?�璺虹灱绾惧ジ鏌ｅΟ铏癸紞濠�?呮暬閺岋紕浠﹂崜褉妲堥梺浼欑稻缁诲牓宕�?濡炪倖甯掔€氼剛澹曠紒妯肩闁瑰瓨鐟ラ悘顏堟倵濮橆剚鍤囬柡宀嬬秮瀵剟宕归鏂ゆ�??閿熶粙姊虹紒妯诲蔼闁稿海鏁诲濠氭晲婢跺﹥顥濋梺鍦圭€涒晠宕曢幘缁樺€垫繛鎴炵懅缁犳绱掓潏銊ユ诞闁诡喗鐟╅�?�妤呭焵椤掑嫬绀夐柕鍫濐槹閻撴洘鎱ㄥ鍡�?⒒闁稿孩姊归〃銉╂�?�閼碱剙鈪垫繝纰樺墲閹倹淇婇柨瀣劅闁靛繆妲呭Λ鍐⒑缁洘鏉归柛�?�尭椤啴濡堕崱妤冪懆闁诲孩鍑归崣鍐ㄧ�?????妞ゅ繋鐒﹂敓锟�?闂備胶绮摫鐟滄澘鍟撮�?�鏃堝Χ婢跺鍘�???妞ゆ劧绲界喊宥咁渻閵堝骸浜濈紒璇茬墦楠炲啫鈻庨幙鍐╂櫌闂�?€炲苯澧存い銏℃閿燂拷???闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹瑩寮堕崹顕呭殭闂傚�?�鍊搁崐鐑芥倿閿曞�?�绠栭柛顐ｆ�?绾炬寧绻濇繝鍌滃閿燂拷?閸愨斂浜滈煫鍥ㄦ尵婢ь澁鎷�??閿熻姤娲樼划�?勫煘閹达附鏅柛鏇ㄥ亗閺夘參姊虹粙鍖℃敾闁搞劌鐏濋悾鐑藉即閵忊€虫濡炪倖甯婄粈浣规償婵犲洦鈷戦柛鎾村絻娴滄繄绱掔拠鑼㈡い顓炴喘�?�粙濡歌椤旀洟鎮楅悷鏉款棌闁哥姵娲滈懞閬嶅礂缁楄桨绨婚梺闈涱槶閸庤櫕鏅跺☉姘辩＜缂備焦顭囧ú�?�橆殽閻愬樊鍎旈柟顔界懅閹瑰嫭绗熼娑辨（婵犵绱曢崑鎴�?磹瑜忓濠冪鐎ｎ亞顔愬銈嗗姧缁犳垿鎮￠敓锟�?閺岀喐娼忛崜褏鏆犻梺缁樻惈缁绘繈寮诲☉銏犵労闁告劧缂氬▽顏嗙磽娴ｉ潧濡块柛妯犲浄鎷�?閿熶粙宕�?鍢壯囨煕閹扳晛濡兼い顒€鐗撳娲箰鎼淬垹顦╂繛�?�樼矤娴滄繃绌�????婵☆垵鍋愰幊婵嬫⒑闁偛鑻晶顔姐亜閺囶亞绉い銏�?�哺閿燂�??閿燂�???闁伙絿鍏�?幃鈩冩償濡粯鏉搁梺璇插嚱缂嶅棙绂嶅┑�?�辈妞ゅ繐鐗婇埛鎺楁煕鐏炲墽鎳呮い锔肩畵閺�?喓鍠婇崡鐐扮盎闁绘挶鍊濋弻鏇熺箾閻愵剚鐝旈梺姹囧€ら崳锝夊蓟濞戞粠妲煎銈冨妼閹虫劗鍒掓繝姘兼晬婵炴垶姘ㄩ鏇㈡倵閻熸澘顥忛柛鐘虫礈閼鸿鲸绺介崨濠勫幗闂佽宕樺▔娑㈠几濞戙垺鐓涢敓锟�?鐎ｎ剙鍩岄柧浼欑秮閺屾稑鈹戦崱妤婁患缂備焦顨忛崣鍐潖濞差亝鍋傞幖绮规濡本绻涚€涙鐭ゅù婊庝簻椤曪絿鎷犲ù瀣潔闂�?潧绻掓慨鐢杆夊┑瀣厽闁绘ê鍘栭懜顏堟煕閺傚潡鍙勭€规洘绻堥�?�娑㈡�??????婵犵數鍋涢悧鍡涙倶濠靛鍑犻柣鏂垮悑閻撴瑦銇勯弮鍌氬付闁逞屽墮濞硷繝骞冩导鎼晩闂佹鍨版禍楣冩煥濠靛棝顎楅柡�?�枛閺岋繝宕ㄩ鍓х厜闂佸搫鐭夌紞渚€寮幇鏉垮窛闁哄顑欐导鍐�?繆閵堝洤啸闁稿鍋ゅ畷婵嗏枎韫囷絾缍庨梺鎯х箺椤�?鎷�?閿熻姤宀搁弻鐔虹磼濡櫣鐟ㄥ┑顕嗙稻閸旀妲愰幘璇茬＜婵ɑ鐦烽姀鈥茬箚妞ゆ劧绲块幊鍛磼椤旂⒈鍎忔い鎾冲悑�?�板嫭绻濋崶褎鏆梻鍌欑閹碱偄煤閵娾晛绐楅幖娣�?灮椤╁弶淇婇妶鍛櫤闁抽攱鍨圭槐鎺炴�??閿熺瓔鍘界涵鍓佺磼閻樺啿鈻曢柡灞界Т閻ｏ繝骞嶉纰辨毇闂備礁纾划顖炲箰閼姐�?�鐭夐柟鐑樻煛閸嬫捇鏁愭惔鈥茬敖闂佸憡眉缁瑥顫忔ウ瑁や汗闁圭儤鍨抽崰濠囨⒑閹肩偛濡洪柛妤佸▕楠炲棝宕橀鑺ュ劒闂侀潻�?�岄崢楣冩晬濠婂牊鈷戠紓浣光棨椤忓嫀鐔哥�?閸ャ劌浜楁繝闈涘€搁幉锟犳偂閿燂�???閸忓浜鹃梺閫炲苯澧寸€规洑鍗冲浠嬵敇濠ф儳浜惧ù锝囩《閺嬪酣鏌熼悙顒佺稇濞寸姴銈搁幃妤呭礂婢跺﹣澹曢梻渚婃嫹?閿熻棄鑻晶鎾煙椤旂懓澧茬€垫澘�?�伴獮鍥敇濞戞瑥顏归梻鍌欐祰�?�曠敻宕伴幇顓犵彾闁糕剝绋掗弲顒婃嫹?閿熷鍎遍ˇ浼存偂閺囥垺鍊甸柨婵嗗暙婵″ジ鏌嶈閸撴岸鎮уΔ鍐煔閺夊牄鍔庨敓锟�?闂佹悶鍎崝�?勫焵閿燂�??椤兘寮婚妶澶婄畳闁圭儤鍨垫慨鏇炩攽閻愬弶鍣规俊顐ｇ〒濡叉劙骞樼€涙ê顎撻梺闈╁瘜閸樼ǹ危閸繍娓婚柕鍫濇閻忋儵鎮�?顐㈠祮閿燂�??????妞ゆ棁妫�??婵犳碍鐓犻柟顓熷笒閸�?鏌熷畡閭︾吋婵﹨娅ｇ划娆撳箰鎼淬垺�?�抽梻浣虹帛濡繘宕滈悢鑲╁祦闊洦绋掗弲鎼佹煥???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鎹愵嚙閻ょ偓銇勯幇鈺嬫�??閿熶粙宕瑰┑瀣厱妞ゆ劗濮撮崝婊堟煛閸涱喗鍊愰柡灞诲姂閹�?�宕掑☉姗嗕�??婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；闁绘劗鍎ら崑�?�煟濡崵�?介柍褜鍏涚欢姘嚕閹绢喖顫呴柍鈺佸暞椤忕喖姊绘担鑺ョ《闁革綇绠撻敓锟�?????缂傚倸鍊烽懗鍫曞磻閹捐纾跨€规洖娲ㄧ粈濠傗攽閻樺弶鎼愰柦鍐枑缁绘盯骞嬪▎蹇曞姶闂佽桨�?�?崯鎾蓟閵娿儮鏀介柛鈩冿供濡�?�顪冮妶蹇氱闁稿骸纾Σ鎰板箳濡や緤鎷�?閿熻姤銇勯幒鍡椾壕闂佸憡鏌ｉ崐妤冩閹炬剚鍚嬮柛婊冨暢閸氼偊鎮楀▓鍨灈妞ゎ厾鍏樺畷瑙勩偅閸愩劎鐤€婵炶揪绲介幉锟犲磹椤栫偞鈷掑ù锝呮啞閸熺偛銆掑顓ф疁鐎规洖缍婇、娑樷堪閸愩劎浜伴梻浣圭湽閸ㄥ綊骞夐敓鐘冲亗闁绘梻鍘х粻瑙勭箾閿濆骸澧�?柣蹇ｅ櫍閺屾盯鎮㈤崫銉ュ绩闂佸搫琚崝鎴�?箖閵堝纾兼繛鎴烇供閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚缁犵偤鎸婇悢鍏肩厪閿燂拷?????闂佺粯鎸婚惄顖炲箖閿燂拷?閹瑩骞撻幒鍡樺瘱闂備線娼уΛ娆戞暜閹烘绠掗梻浣虹帛閻熴儵骞婇幇鐗堝仼闁汇垻顣介崑鎾舵喆閸曨剛顦ㄧ紓渚囧枛缁绘ǹ妫熷銈嗘⒐閸ㄦ繄鎹㈤崱娑欑厵缂備焦锚缁椦冾熆瑜庡ú姗€濡甸崟顖ｆ晜闁告洦鍋呭▓缁樼節閿燂�???瀹曞洤鐓熼悗瑙勬磸閸斿酣鍩€椤掑倹鏆�??濠碉紕鍋樼划娆忣潖缂佹ɑ濯撮柣鎴灻▓�?勬⒑閹肩儑鎷�??閿熶粙鎮ч悩鑽ゅ祦闊洦绋掗弲鎼佹�???
    
        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺妫冨畷鍗炩枎閹搭垳搴婄紓鍌氬€搁崐鐑芥�?�閿曞偊鎷�?閿熶粙宕堕�?�鈩冩そ楠炴﹢顢欓悾灞藉箥闁诲氦顫夊ú鏍洪妶澶婄厺闁割偆鍠嗘禍婊堟煏韫囧﹥顫婇敓锟�?????闁哄洨鍠庣粭鎺撱亜椤愶絿绠栨い顐ｅ灴瀵€燁槺閺夆晜锕㈠濠氬磼閿燂�???閹间礁纾归柣鎴ｅГ閸ゅ嫰鏌ら崫銉︽毄濞寸姵纰嶆穱濠囨�??????闂佹悶鍔庨弫璇茬暦椤栫偛绾ч柟瀵稿У濞堥箖姊洪崫鍕偍闁搞劍妞藉畷鎴�?Ω瑜忛敓锟�?????妞ゆ挾鍋涙慨鐑芥⒑绾懎袚婵炶尙鍠庨～蹇撁洪鍕唶闁硅壈鎻徊鍧楁偩闂堟侗娓婚柕鍫濈箰閻︽粓鏌涢妸銉у煟闁轰焦鍔欓幃娆撳传閸曨偆鐛╅梺璇插缁嬫帡鈥﹂崶顒€鍌ㄩ柟鍓х帛閻撴稑顭跨捄楦垮濞寸媴绠戦埞鎴︻敍濞嗘垹鐓撻悗瑙勬礃椤ㄥ牊绂掗敃鍌涘剹妞ゆ劑鍨荤粔娲煙椤旂懓澧查柟顖涙閿燂拷?闁绘ê纾禍宄扳攽閻樻剚鍟忛柛鐘崇墵閺佸啴濡烽妷顔藉瘜闂佽姤锚椤﹂亶寮抽敂濮愪簻闁规澘澧庨悾閬嶅船椤栫偞鈷戦梻鍫熶緱濡插綊鏌涢弬鐐叉噹缁躲倕螖閿濆懎鏆欏鍛存⒑閸涘﹥澶勯柛銊у閸庮偊姊绘担鐟邦嚋婵炴彃绉瑰畷鎴﹀箻閺傘儲鏂€濡炪倖妫�?崑鎰墡婵＄偑鍊戦崝濠囧磿閻㈢ǹ绠栨繛鍡樻尰閸ゆ垶銇勯幒鎴濅簽闁哥喎顑夊缁樻媴閼恒儻鎷�?閿熶粙鏌ｉ幒鐐电暤妤犵偞鍨垮畷鍫曨敆?闁哄绶氶弻鐔煎礈瑜忕敮娑㈡煛閸涱喗鍊愰柡灞诲姂閹倝宕掑☉姗嗕�???闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩冾殔琚濋梻浣告啞閹稿爼宕濋幋锔惧祦闊洦绋掗弲鎼佹煥???闂傚倸鍊峰ù鍥р枖閺囥垹绐楃€广儱娲ら崹婵囩箾閸℃绂嬫繛鍏肩墬缁绘稑顔忛鑽ゅ嚬闂佸搫鎳忛幃鍌炲蓟閵娾晜鍋嗛柛灞剧☉閿燂拷??缂傚倸鍊搁崐椋庣矆閿燂拷?钘濇い鏍剱閺佸銇勯幘璺盒㈤柛銊︾箓閳规垿鎮╅崘鎻掓瘓闂佽桨绀佺粔褰掑蓟閿濆绠涙い鎺戭槸濞堝爼姊洪崨濞楃懓螞閸曨垰鐓�?柟杈剧畱閻擄繝鏌涢埄鍐炬畼濞寸媭鍘奸—鍐Χ閸℃浠搁梺鑽ゅ暱閺呮盯鎮鹃悜鑺ヮ棃婵炴垶甯楅悗濠氭⒑閻熼偊鍤熷┑顔惧厴閺佸秴饪伴崼鐔叉嫼缂傚倷鐒﹂敃鈺呮倿娴犲鐓涘ù锝呮啞閹叉悂鏌℃笟鍥ф灈闁宠棄顦甸敓锟�??闁挎稑�?�敮楣冩⒒娴ｈ鍋犻柛搴㈢矒�?�曟﹢宕ｉ妷褏锛為梻浣筋嚙鐎涒晠顢欓弽顓為棷??鐎规洘濞婇弫鎰板川椤栨稒顔曢梻浣稿閸嬪懎煤瀹ュ鐒垫い鎺嶈兌婢у灚銇勯姀锛勬噰闁瑰磭鍋ゆ俊鐑藉�?????缂傚倸鍊搁崐鐑芥嚄閸撲礁鍨濇い鏍仦閸庡孩銇勯弽銊︾殤闁哄棴绠撻弻鏇熺箾閻愵剚鐝﹂梺杞扮閸熸挳寮婚弴锛勭杸闁挎繂妫涚粣鏃傜磽娴ｄ粙鍝洪柣鐕傚閹广垹鈹戦崱蹇旂亖闂佸壊鐓堥崰妤呮�?�閸儲鈷戦柟绋垮绾炬悂鏌涙惔銊ゆ�????闂佸憡鍔﹂崰妤嬫�??閿熺晫濮撮�?�璺ㄦ崉閻戞ɑ鎷卞┑鐐茬墛閸庢娊鈥旈崘顔嘉ч柛鈩冾殔琛肩紓鍌欒兌婵敻宕归崷顓炲灊闁割偀鎳囬崑鎾绘晲鎼粹€茬按婵炲瓨绮嶇划鎾诲蓟閻斿吋鐒介敓锟�??闁哄鐩弻鈽呮�??閿熺瓔浜妤呮婢跺绡€濠电姴鍊绘晶銏ゆ煟閿濆棙銇濋柡宀嬬磿娴狅箓宕滆閸掓稑顪冮妶鍐ㄧ仾婵炶尙鍠栧顐�?箛閺夊灝鑰垮┑鐐叉钃辩悮锝囩磽閸屾熬鎷�??閿熶粙鎳楅崼鏇炵；闁规崘顕х壕鍖℃�??閿熻姤娲栧ú銊х矆婵犲�?�鏀介柣妯哄级閹兼劙鏌﹂崘顏勬灈闁哄苯绉归敓锟�???濠⒀屽灦閺屾稑顫濋澶婂壎闂佸搫鏈粙鎴�?煡婢舵劕纭€闁绘劕鍚€閹撮绱撻崒娆戣窗闁哥姵宀稿顐ｇ�?濮橆剝鎽曢梺鎸庣箓濡瑩宕曢悢鍏肩厪闊洤顑呴悘鈺呮煛閸☆厾绡€婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘�?閿燂�??????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑掳鍊曢崯顐﹀垂濠靛棌�?介柣妯虹枃婢规绱掗悪娆忔搐缁犲綊鎮�?☉娅虫垹浜告导�?�樼厸闁稿本顨呮禍楣冩⒒閸屾熬鎷�??閿熶粙鎳楅崜浣稿灊妞ゆ牜鍋為弲顏堟煟鎼淬埄鍟忛柛鐘崇墵閹儲绺介崫銉ョウ闂佸搫绋�?崢鑲╃不濞戙垺鐓�???闁绘绻樺畷銏ゅ�?閻愨晜鏂€闁圭儤濞婂畷鎰板箻閸撲胶鐒兼繛鎾村焹閸嬫捇鏌涢埞鍨伈鐎殿喗鎸抽敓锟�?闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣枛�?�曟垿骞�?崜浣虹劶婵犮垼娉涢惉鑲╁婵傚憡鐓熸俊顖濇閿涘秹鏌嶉娑欑缂佽鲸甯炵槐鎺懳熼懖鈺冩澖闁诲氦顫夊ú妯兼暜閹烘缍栨繝闈涱儐閺呮煡鏌涢埄鍐炬畼鐟滅増鍎抽埞鎴︽偐閸偅姣勬繝娈垮枤閸忔ê顕ｉ锕€绠瑰ù锝呮憸閿涙稑鈹戦悙鏉戠仧闁搞劌�?辩划濠氭偐绾版ê浜鹃柛蹇擃槸娴滈箖姊洪崨濠冨闁稿�?�伴幃妤咁敇閵忊檧鎷洪梺鍏间航閸庡秹顢旈崺璺烘喘閹稿﹥寰勫Ο鐓庡Ш闂備礁鎼粙渚€宕㈡禒瀣亗闁挎繂顦遍崣鎾绘煕閵夛絽濡奸柛銈庡墯缁绘盯宕楅悡搴☆潕闂侀€炲苯澧叉い顐㈩槸鐓ら柡宥庡帞閸ヮ剚鍋ㄧ紒�?�劵閹芥洟姊洪崫鍕�?窛闁哥姵鎸剧划缁樸偅閸愨晝鍘卞銈庡幗閸ㄧ敻寮稿☉妯锋斀妞ゆ棁濮ょ粈瀣叏婵犲懏顏犵紒杈ㄥ笒铻ｉ柤娴嬫櫇缁愭姊绘担瑙勫仩闁告柨绻愯灋闁告洦鍨界紞鏍叓閸ャ劎鈯曢柟顖滃仱閹嘲鈻庤箛鎿冧患缂佸墽铏庨崹璺侯潖濞差亝顥堟繛娣�?妼缂嶅﹤鐣烽弴銏犺摕闁靛�?绠戞禒褔姊洪棃娑氱疄闁稿﹥鐗犻崺娑㈠箣閿旂晫鍘介梺缁樻煥閹诧紕娆㈤崣澶岀闁割偅纰嶅▍濠囨煛鐏炶濮傞柟顔哄€濆畷鎺戔槈濮楀棔绱�???
        .ex_bpu_is_bj(ex_is_bj),
        .ex_pc1(ex_pc1),
        .ex_pc2(ex_pc2),
        .ex_valid(ex_valid),
        .ex_bpu_taken_or_not_actual(ex_real_taken),
        .ex_bpu_branch_actual_addr1(ex_real_addr1),  
        .ex_bpu_branch_actual_addr2(ex_real_addr2),
        .ex_bpu_branch_pred_addr1(ex_pred_addr1),
        .ex_bpu_branch_pred_addr2(ex_pred_addr2),
        .get_data_req_o(get_data_req),
        .csr_dmw0(csr_dmw0),
        .csr_dmw1(csr_dmw1),
        .csr_da(csr_da),
        .csr_pg(csr_pg),
        .csr_plv(csr_plv),

/*******************************
        .tlbidx(),
        .tlbehi(),
        .tlbelo0(),
        .tlbelo1(),
        .tlbelo1(),
        .asid(),
        .ecode(),

        .csr_datf(),
        .csr_datm(),
***********************************/

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚缁犵偤鎸婇悢鍏肩厪閿燂拷?????闂佺粯鎸婚惄顖炲箖閿燂拷?閹瑩骞撻幒鍡樺瘱闂備線娼уΛ娆戞暜閹烘绠掗梻浣虹帛閻熴儵骞婇幇鐗堝仼闁汇垻顣介崑鎾舵喆閸曨剛顦ㄧ紓渚囧枛缁绘ǹ妫熷銈嗘⒐閸ㄦ繄鎹㈤崱娑欑厵缂備焦锚缁椦冾熆瑜庡ú姗€濡甸崟顖ｆ晜闁告洦鍋呭▓缁樼節閿燂�???瀹曞洤鐓熼悗瑙勬磸閸斿酣鍩€椤掑倹鏆�??濠碉紕鍋樼划娆忣潖缂佹ɑ濯撮柣鎴灻▓�?勬⒑閹肩儑鎷�??閿熶粙鎮ч悩鑽ゅ祦闊洦绋掗弲鎼佹�??? dcache 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幏鐘绘嚑椤掑偆鍞洪梻浣呵归敓锟�???濡炪們鍨烘穱娲�?�囪ぐ鎺撶厱闁宠鍎虫禍鐐繆閻愵亷鎷�?閿熺晫鏁繝鍕偨闁炽儲鏋奸弸鏃€绻濇繝鍌滃�?闁绘挶鍎甸弻锝夊�??????????濠电姷顣槐鏇㈠磻閹达箑纾归柡宥庡亝閺嗘粌鈹戦悩鍙夊闁搞�?��?�伴弻娑㈩敃閿濆棛顦ラ梺缁樻尨閸嬫捇姊绘担鍛婃儓婵炲眰鍨藉畷褰掓惞閸忓浜炬慨姗嗗墯閸ゅ洦鎱ㄦ繝鍐┿仢妞ゃ垺顨婇敓锟�??妞ゆ帒鍊婚惌鎾绘煟閵忕姵鍟為柛�?�€块弻锝夊棘閸喗鍊梺缁樻尭缁绘劙鍩為幋锔藉亹闁肩⒈鍓涢濠囨⒑娴兼瑧绉ù婊冪埣�?�鏁愰崼銏㈡澑闂佸搫鍟犻崑鎾绘�?�韫囥儳鐣甸柡宀嬫嫹?閿熺晫鏆嗛柍褜鍓熷畷浼村�?????濠电偛妫欓崹鍫曞窗閸℃稒鐓欓柣鎴灻悘锕傛偣閹板墎纾跨紒杈ㄥ浮椤㈡瑥鈻庨幆褎顔勯梻浣哥枃濡嫰藝椤栫儑缍栨繝闈涱儐閺呮煡鏌�???妞ゃ儲宀稿缁樻媴閻熼偊鍤嬬紓浣筋嚙閸婂鎳為柆宥嗗殐闁冲搫瀚皬缂傚�?�鍊烽悞锕佸綘婵炲瓨绮嶇划宥夊Φ閸曨垰绠涢柍杞拌兌娴犻箖姊洪悷鏉挎倯闁告梹鐟╅獮妤呭醇閺囩偛鍞ㄥ銈嗘尵閸犳捇宕㈤挊澶嗘斀妞ゆ柨顫曟禒婊堟煕鐎ｎ偅灏扮紒缁樼⊕閹峰懘宕�?幓鎺濅紑濡炪倐鏅犻弨杈╂崲濠靛洨绡€闁稿本绋戝▍褏绱掗悙顒€�?冮柛瀣姉濡叉劙骞樼€涙ê顎撻梺璋庡惓褰掑矗閺囥垺鈷戦柛蹇曞帶椤庢粍绻涙径瀣�???濡炪倖甯婄欢锟犲疮韫囨稒鐓曢柨婵嗛�?�濞呭稄鎷�?閿熻姤娲�?崹鍓佹崲濠靛鐐婄憸搴ㄦ倵椤掑嫭鈷戦柣鐔告緲閳锋梻绱掗鍛仸鐎殿喗鐓￠獮鏍ㄦ媴閸︻厼寮抽梻浣虹帛濞叉牠宕�???????
        .ren_o(backend_dcache_ren),
        .wstrb_o(backend_dcache_wen),
        .writen_o(backend_dcache_writen),
        .virtual_addr_o(backend_dcache_addr),
        .wdata_o(backend_dcache_write_data),

        // dcache 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倸鍊风欢姘跺焵椤掑�?�浠滈柤娲诲灡閺呰鎷�?閿熺晫纭堕崑鎾舵喆閸曨剛锛涢梺鍛婎殔閸熷潡顢氶敐鍡欘浄閻庯絽鐏氶弲锝夋⒑缂佹〒鍦焊濞嗘挸围闁挎洖鍊归埛鎺懨归敐鍛暈闁诡垰鐗忕槐鎺炴嫹?閿熻В鏅濈粣鏃撴嫹?閿熻姤娲╃徊楣冨箚閺冨牆惟閿燂拷?????闂傚倷鐒﹂幃鍫曞磿椤栫偛�?夐幖杈剧到婵剟鏌嶈閸撶喎顫忔繝姘＜婵ê宕敓锟�??缂傚倷绀�?鍡涘箰婵犳艾鐤鹃悹楦裤€€濡插牓鏌曡箛銉х？闁告ɑ鎮傚娲川婵犱胶绻�?梺鍛娒妶鎼佺嵁閸愵喖绠ｆ繝鈧灩闁帮絽鐣烽幆閭︽�?�闂傚⿴鍓﹂崜鐔煎蓟閻旂⒈鏁婇柣锝呮湰閸ｆ澘顪冮妶鍐ㄧ仾婵☆偄鍟悾鐑芥偄閻撳宫鈺呮煏婢跺牞鎷�?閿熶粙藟濮樿埖鐓熼柣鏂挎憸閻﹦绱掔紒妯虹瑨閸楅亶鏌熼幍顔碱�????闂備礁鎲＄换鍌︽�??閿熺瓔鍓熼幊鎾诲垂椤旇鏂€闂佺粯鍔栧娆撴倶閿曞�?�鐓ラ柡鍥悘鈺呮懚閻愮儤鐓熼柟杈剧到琚氶梺鎶芥敱閸ㄥ潡寮婚悢铏圭煓闁圭ǹ�?�╁畷宕囩磽娴ｅ搫校闁圭ǹ顭锋俊鐢稿礋椤栨稒娅囬敓锟�????闁伙絿鍏�?、妤呭礋閿燂�??娴犲ジ姊哄Ч鍥х仼闁硅绻濆鏌ュ箹娴ｅ湱鍙嗛梺缁樻�?閿燂�?????闂傚倸鍊烽懗鍓佸垝椤栫偛绠归柍鍝勬噹绾捐鈹戦悩璇ф嫹?閿熶粙寮抽敃鍌涚厱妞ゆ劧绲鹃敓锟�??闁诡垳鍠栭幃宄扳堪閸愮偓效闂�?€涚┒閸�?垵鐣烽崼鏇ㄦ晢濞达絽寮剁€氳偐绱撻崒娆戭槮妞ゆ垵鎳愭禍鎼佸川椤撗冩櫊闂侀潧顧€鐠愮喐绂嶅⿰鍕�?簻闁规崘娉涘瓭闂佸憡锚椤曨參鍩€椤掍緡鍟忛柛鐘崇墵閳ワ箓鏌ㄧ€ｂ晝绠氶梺鍏兼倐濞佳呮閻愭祴�?介柣妯诲絻椤忣偊鏌￠崱鎰伈婵﹦绮幏鍛村川婵犲懐顢呴梻浣呵圭花娲磹濠靛棛鏆︾憸鐗堝笒閸ㄥ�?�銇勯幇鍓佸埌鐎殿喖娼�?�娲传閸曨剙绐涢梺绋款儐閸旀瑥顕ｉ妸锔绢浄閻庯綆鍋嗛崢浠嬫⒑瑜版帒浜伴柛鎾寸懅閻ヮ亣顦归柡灞剧洴閺佹劙宕惰楠炲姊洪崫鍕拱闁烩晩鍨辨穱濠囧箹娴ｈ倽鈺呮煥閺冨倻甯涙い銉ヮ槹娣囧﹪鎮�????闂佺ǹ顑呯€氼噣骞戦姀銈呯�?妞ゆ梻鍘ч悿鎯р攽閿涘嫬浜�???缂備胶绮崝娆撶嵁婵犲啯鍎熼柕蹇嬪焺濞茬ǹ鈹戞幊閸婃洟骞婅箛娑欏亗婵炲棙鎸婚悡鐘绘煕閿旇骞栨い锝堝亹閹叉悂骞庢繝鍌涘櫧缁炬儳銈搁弻锛勪沪鐠囨彃濮㈤梺浼欑悼閸庛�?�銆冮妷鈺傚€烽敓锟�?????闂備浇顕栭崰鎺楀礈濠靛绠氶柡鍌濐嚦閻旇櫣纾兼俊顖滅帛缁额偅绻濈喊澶�?？闁稿鍨垮畷鎰板冀椤剚绋掔粭鐔煎焵椤掑嫭鏅查柣鎰�?棘閺冨牆鐒垫い鎺戝閸嬫垵霉閸忓吋缍戦梺鍗炴处缁绘繈妫冨☉姘拡濠德ゅ皺閸忔ê顫忓ú顏呭仭闁哄瀵ч崐顖炴⒑娴兼瑧绉靛ù婊庝簻閻ｉ鎲撮崟顓犵槇濠殿喗菧閸庮噣宕戦幘璇插窛闁哄鍨奸幗鏇㈡⒑闂堟侗妾у┑鈥虫喘瀹曘垽鎮介崨濞炬嫽闂佺ǹ鏈懝楣冨焵椤掍焦鍊愭い銏″哺椤㈡﹢鍩楅崫鍕枠闁轰礁鍟村畷鎺戭潩鏉堚晜姣庨梻鍌欒兌缁垶寮婚妸鈺佽Е閻庯綆鍠栭悡鏇㈡煙鏉堥箖妾�?柛濠勬暬閺屾盯鏁傜拠鎻掔闁哄稄绻濆娲濞戞瑯妫為梺鍝ュ枑閹稿啿顕ｆ繝姘у璺猴功椤︺劑姊洪懖鈹炬嫛闁告挻鐟╅幃锟犳偄婵傚瀵岄梺闈涚墕閸燁偊鎮�?鍫熺厽闁绘柨寮跺▍鍛存煟閿濆洤鍘寸€规洩绻濋幃娆撳煛閸屻�?�缍屽┑鐘垫暩閸嬫稑螞濞嗘挸鍨傞梻鍫熶緱閸ゆ洟鏌熼幆鏉啃撻柍閿嬪笒闇夐柨婵嗙墛椤忕娀鎮介娑氣姇缂佺粯鐩畷锝嗗緞鐏炶В鎷伴柣搴ゎ潐濞叉﹢宕濆▎鎾崇畾闁稿瞼鍋涘婵嗏攽閻樻彃浜�???闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柟鐗堟緲閸戠姴鈹戦悩瀹犲缂佺媭鍨堕弻銊╂偆閸屾稑顏�???
        .rdata_i(dcache_rdata),
        .rdata_valid_i(dcache_backend_rdata_valid),
        .dcache_pause_i(~dcache_ready),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠囧极瀹ュ拋鍚嬮柛鈩冩礈缁犳岸姊洪崨濠勬噧妞わ富鍨遍幈銊ヮ吋閸�?晜顔旈梺缁樺姈濞兼瑥霉閿燂拷??濞堝灝娅�?柛鎾跺枛楠炲啫鈻庨幙鍐╂櫌闂�?€炲苯澧柛鎺戯躬楠炲秹顢欓崜褝绱抽梻浣呵归張顒勬偡瑜斿畷婵嗩吋閸モ晝锛滈柣搴秵閸嬪嫰鎮樼€涙ǜ浜滈柕蹇ョ磿婢х鎷�?閿熻姤娲樼敮锟犲箖濞嗘挻鍤戞い鎺戯功楠炪垽姊婚崒娆愮グ妞ゎ偄顦敓锟�????妞ゃ垺淇洪ˇ褰掓煙椤旀儳浠遍柟顔荤矙�?�曘劍绻濋崟顐㈢闂傚�?�鑳剁划顖氼潖绾懌浜归柛鎰ㄦ櫇椤╄尙绱掔捄鐑樺枠婵﹤顭峰畷鎺戭潩椤戣棄浜鹃柟闂寸绾惧綊鏌熼梻�?�割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繑鎸抽弻锛勪沪閸撗€妲堥梺�?�狀潐閸ㄥ灝鐣烽崡鐐嶆梹绻濇担铏癸紳闂傚倷娴囬褝鎷�??閿熻В鏅涢～婵嬪Ω閿旇姤鐝峰┑掳鍊曢幊搴㈩攰闂備礁鎲″ú锕傚垂闁秴鐤炬繝濠傜墛閸嬶綁鏌涢妷顔荤盎闁汇劌鎼湁闁绘ǹ娅曠亸锔芥叏婵犲懏顏犻柟椋庡█閹崇娀顢楅崒銈呮暪濠碉紕鍋戦崐鏍垂閻㈡潌鍥敍閻戝洨绋忛棅顐㈡处閹峰煤椤忓秵鏅滈梺鍛婃处娴滅偤鎮欐繝鍥ㄢ拻濞达絽鎲￠崯鐐寸箾鐠囇呯暤鐎规洘鍨垮畷銊╊敇濞戞瑧浜栨俊鐐€栭幐鍫曞垂濞差亜鐓曢柟瀵稿Х绾捐棄霉閿濆洦顏熷�?�姘⊕缁绘盯宕奸悢鍓叉闂佸搫琚崝鎴濐嚕閹绢喖惟闁靛牆娲ㄥ▔鍧楁⒒娴ｉ涓茬紒鎻掓健閿燂�????閿燂�??????妞ゆ棁妫勬禍鐟邦渻閵堝棗濮﹂敓锟�???婵犮垼顫夊ú鐔奉潖濞差亜绠伴幖杈剧悼閻ｅ灚淇婇妶鍥㈤柟璇х磿缁顓兼径�?�舵�??閿熶粙鏌ｉ姀銏℃毄闁挎稒绮撳铏圭磼??閻庤娲滈弫濠氬箖閹灐娲敂閸涱垰骞�???闁�?�屽墴閿燂拷?妞ゆ帒�?�梻顖炴煥閺囩儑鎷�??閿熺晫绮婚鐐寸叆閿燂拷?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵愭Т闁�?�屽墾缁犳挸鐣烽崼鏇ㄦ晢闁�?�屽墰缁鎮╃紒妯煎幈闂侀€涘嵆濞佳囧几閻斿吋鐓熼柟鎹愭硾閺嬫盯鏌ｉ幙鍐ㄤ喊鐎规洝鍩栭ˇ鐗堟償閳藉棗娈奸梻鍌氬€风欢锟犲矗鎼淬劌鍨傞柛顐ｆ礀閽冪喖鏌嶉妷銉э紞闁哄棗妫濋幃妤呮晲鎼粹€愁潾闂佷紮绠戦悧鎾诲箖濡ゅ啯鍠嗛柛鏇ㄥ墰閿涙﹢姊洪崨濠冣拹闁搞劌娼℃俊�?�樻媴缁洘鐎婚梺鍦亾濞兼瑩鎯傞崟顒傜瘈闁靛骏绲剧涵鐐繆椤愶綆娈曠紒鍌氱У閵堬綁宕�?埡鍐ㄥ箥闂備浇顫夐鏍窗閺嶎叏鎷�?閿熻姤绺介崨濠勫幗闂佽鍎抽顓灻洪幘顔界厵妞ゆ梹鏋婚懓鍧楁煙椤旂晫鎳勯柨娑欏姇閳规垿宕卞鍡楁暢濠电姷鏁告慨鐢割敊閺嶎厼绐楅柡宥庡幖绾惧綊鏌涜椤ㄥ懘鎷戦悢鍏肩厽闁哄啫鍊甸幏锟犳煛娴ｉ潻韬柡宀嬬到椤繈顢楅崒娑欏枛闂佽瀛╅敓锟�?????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牗绋戞禒濂告⒑缂佹ê鐏辨俊顐㈠缁骞庨懞銉у幍闁诲孩绋掕摫闁抽攱鍔栭妵鍕敃閵忊懣銏ゆ煃鐟欏嫬鐏存い銏＄懅缁鎷�??閿熺瓔鍋嗛弳銉︾�?绾版ɑ顫婇柛�?�噹铻為柛鎰靛枛閺嬩線鏌熼崜褏甯涢柡鍛�?�閺屻劑鎮ら崒娑橆伓?8濠电姷鏁告慨鐑藉极閸涘﹥鍙忛柣鎴ｆ閺嬩線鏌涘☉姗堟敾闁告瑥绻橀弻锝夊箣閿濆棭妫勯梺鍝勵儎缁舵岸寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ゆい顓犲厴�?�鏁愰崨鍌滃枎閳诲酣骞嗚椤斿嫮绱撻崒娆掑厡濠殿喗鎸抽幃妯侯潩鐠轰綍锕傛煕閺囥劌鏋�??闂備礁婀遍崑鎾诲箚鐏炶娇娑㈡倷閻㈢數锛濇繛杈剧悼閺咁偊宕奸鍫熺厱濠电姴鍟扮粻鐑囨嫹?閿熺瓔鍠栭�?�鐑藉极閹邦厼绶為悗锝庡亝閻濇娊姊绘担鍛婂暈濞撴碍顨婂畷褰掓惞椤愩埄鍤ら梺鎼炲労閸撴岸鍩涢幋鐐电闁煎ジ顤傞崵娆愵殽閻愭惌娈滈柡�?€鍠栭獮鏍ㄦ媴閾忚姣囨俊銈囧Х閸嬫盯藝閻㈠摜宓侀柡宥冨妽婵挳鏌ｉ悢纰辨殥缂傚啯娲熷缁樻媴缁嬫妫岄梺绋款儏閹虫劙骞戦�?銈呯妞ゆ牗绋戞禒顓㈡⒑闂堟单鍫ュ疾濠婂牆鐓曢柟杈鹃檮閻撴洘绻濋棃娑欘棞妞ゅ繑鎸抽弻娑欐償閳╁啯宕崇紓浣介哺鐢繝骞婂⿰鍫燁棃婵炴垶蓱閹虫瑩鏌ｆ惔銏╁晱闁哥姵鐗犻垾锕傛倻閽樺鐣洪梺闈涚箞閸婃牠宕戦崒鐐茬閺夊牆澧界粔鐢告煕閻愯尙绉烘慨濠勭帛缁楃喖鍩€椤掑嫬鐒垫い鎺嶈兌閳藉鎷�?閿熻姤鎸稿Λ娆戞崲濞戞瑦濯撮柛鎰絻閺嗗﹪鏌＄€ｎ偅鈷愰柕鍥у楠炴鎹勬潪鐗堢潖闂備浇銆€閸嬫挸霉閻樺樊鍎愰柣鎾冲暣閺岋箑螣娓氼垱效濡炪�?�鍎茬划�?勬箒濠电姴锕ょ€氼喚绮婚悙鐑樼厸閻忕偠顕ф慨鍌︽嫹?閿熺瓔鍠�?娆掔亽閿燂�??????缂佽鲸鐟╅弻锝嗘償閵忊晛鏅遍梺鍝ュУ閿燂拷????閻庣懓�?�伴崑濠囧吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏″殗闁哄矉绲借灒婵炲棙鍎冲▓顓㈡⒑鏉炵増绁版い顐㈩槺閹广垹鈹戠€ｎ偄浠洪梻鍌氱墛缁嬪牓寮搁崨顓涙�?闁绘劖婢樼亸鍐煕韫囨洖孝缂傚秴锕ら悾鐑藉箳閹宠埖甯″畷妤呮嚃閳哄�?�鍨遍梻浣筋嚃閸犳鎮烽埡鍛畺婵犲﹤鍚�?悢鍏肩叆閻庯綆浜舵导鏍⒒閸屾瑦绁扮€规洖鐏氶幈銊╁垂椤愩�?�娲告繛瀵稿Т椤戝懐绮堟径鎰€堕柣鎰礋閹烘鍑犵€广儱顦伴悡娆撴煙濞堝灝鏋涙い锝呫偢閺岋綁骞樼€靛憡鍣伴梺鍝勬湰閻╊垶鐛€ｎ亖鏋庨煫鍥э工娴滈箖鏌″搴�?�簮闁稿鎸搁～婵嬫�?????
        .flush_o(flush_o),
        .pause_o(pause_o),

        .icacop_en(icacop_en),
        .dcacop_en(dcacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),
        
        //debug
        .debug_wb_valid1(debug_wb_valid1),
        .debug_wb_valid2(debug_wb_valid2),
        .debug_pc1(debug_pc1),
        .debug_pc2(debug_pc2),
        .debug_inst1(debug_inst1),
        .debug_inst2(debug_inst2),
        .debug_reg_addr1(debug_reg_addr1),
        .debug_reg_addr2(debug_reg_addr2),
        .debug_wdata1(debug_wdata1),
        .debug_wdata2(debug_wdata2),
        .debug_wb_we1(debug_wb_we1),
        .debug_wb_we2(debug_wb_we2) 
    );

    wire icache_ren_received;
    wire dcache_ren_received;
    wire icache_flush_flag_valid;

    icache u_icache
    (
        .clk(aclk),
        .rst(rst),   
        .flush(flush_o[1]),       
    // Interface to CPU
        .inst_rreq(inst_rreq),  
        .inst_addr1(inst_addr1),   
        .inst_addr2(inst_addr2),  
        .if_pred_addr1(if_pred_addr1),
        .if_pred_addr2(if_pred_addr2),
        .BPU_pred_taken(BPU_pred_taken),

        .icacop_en(icacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),

        .pi_is_exception(pi_is_exception),
        .pi_exception_cause(pi_exception_cause),

        .pred_addr1(pred_addr1_for_buffer),
        .pred_addr2(pred_addr2_for_buffer),
        .pred_taken(pred_taken_for_buffer),
        .inst_valid1(icache_inst_valid1),  
        .inst_valid2(icache_inst_valid2),   
        .inst_out1(icache_inst1),       
        .inst_out2(icache_inst2),
        .valid_out(icache_valid_out),
        .pc1(icache_pc1),
        .pc2(icache_pc2),
        .pc_is_exception_out1(pi_icache_is_exception1),
        .pc_is_exception_out2(pi_icache_is_exception2), 
        .pc_exception_cause_out1(pi_icache_exception_cause1),
        .pc_exception_cause_out2(pi_icache_exception_cause2),
        .pc_suspend(pc_suspend), 
    // Interface to Read Bus
        .dev_rrdy(dev_rrdy_to_cache),       
        .cpu_ren(icache_ren),       
        .cpu_raddr(icache_araddr),      
        .dev_rvalid(icache_rvalid),     
        .dev_rdata(icache_rdata),
        .ren_received(icache_ren_received),
        .flush_flag_valid(icache_flush_flag_valid)   
    );

    wire debug_wb_valid1;
    wire debug_wb_valid2;
    wire [31:0] debug_pc1;
    wire [31:0] debug_pc2;
    wire [31:0] debug_inst1;
    wire [31:0] debug_inst2;
    wire [4:0] debug_reg_addr1;
    wire [4:0] debug_reg_addr2;
    wire [31:0] debug_wdata1;
    wire [31:0] debug_wdata2;
    wire debug_wb_we1;
    wire debug_wb_we2;

    wire [3:0] duncache_wstrb;

    wire cache_axi_write_pre_ready;
    wire duncache_en;

    dcache u_dcache(
        .clk(aclk),
        .rst(rst),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹寸偛顥氶柛娆忔惈閳规垿鎮╅崹顐ｆ瘎婵犳鍠氶崗姗€濡撮崒娑氼浄閻庯綆浜為ˇ顓炩攽閻樼粯娑фい鎴濇噽缁寮介鐔哄幈闁诲繒鍋涙晶浠嬪煟閵壯呯＜閻犲洤寮堕ˉ銏ゆ煛瀹€瀣М妤犵偛顑夐弫鎰板川閸涱喗宕岄柡宀嬬節瀹曘劑顢欓崜褏鍘掔紓鍌欐祰妞存悂骞愭繝姘闁告稑鐡ㄩ崕�?€绱掔€ｎ亞浠㈢憸鏉挎閳规垶骞婇柛濠冾殕閹鳖煉鎷�?閿熻棄鎲″畷鍙変繆椤栨瑨顒熸繛鍏肩墱缁辨挻鎷呴懖鈩冨灦閸掑⿵鎷�?閿熻棄鎽滅壕鍏肩箾閹寸儑渚涢柛搴＄箲缁绘盯宕奸銏犵缂備浇椴搁幐濠氬箯閸涘瓨鎯為柣鐔稿椤愬ジ姊绘担鍛婂暈婵﹤缍婇妴鍐╃�?閸モ晛绁﹂梺纭呮彧缁犳垿锝為崨�?�樼厪闁割偅绻冮崵鍥煕閻愯尙鍩ｆ慨濠冩そ濡啫鈽夋潏銊愩�?�姊虹粙鍨劉濠电偛锕ㄥΛ鐔奉渻閵堝棙纾甸柛�?�尰閹便劍绻濋崨顕呬哗濠电偞鍨归弫璇茬暦閵娾晩鏁婇柛蹇撱偢閺侇亝绻濋悽闈浶ユい锝勭矙閿燂拷?妞ゆ帒鍟悵顏堟煙閸忕厧濮嶉柡宀嬬秮閺佹劙宕堕妸锔界槗闂備浇妗ㄩ悞锕傚箲閸ヮ剙鏋�?柟鍓х帛閺呮悂鏌�???闂傚倸鍊烽懗鍓佸垝椤栫偛绠归柍鍝勬噹绾捐鈹戦悩璇ф嫹?閿熶粙寮抽敃鍌涚厱妞ゆ劧绲鹃敓锟�??闁诡垳鍠栭幃宄扳堪閸愮偓效闂�?€涚┒閸�?垵鐣烽崼鏇ㄦ晢濞达絽寮剁€氳偐绱撻崒娆戭槮妞ゆ垵妫濋、鏍р枎閹惧磭锛熷┑鐐村灦閳笺倝鎮�???闂佸憡娲﹂崢楣冩偪閸曨剛绡€缁炬澘顦辩壕鍧楁煛娴ｇ瓔鍤欓柣锝囧厴閹垻鍠婃潏銊︽珫婵犳鍠楅敃鈺呭礈濞嗘挸鏋�?柕鍫濐槹閳锋帒霉閿濆懏璐￠敓锟�?娴犲鐓曢柕濞垮妽椤ュ銇勯鐐寸┛閿燂�??????闁哄洠鍓濋鐘裁归悪鍛洭闁瑰弶鎸抽弫鎰板幢濡粯绶梻鍌氬€烽懗鍓佸垝椤栫偛绀夋俊顖炴？閻掑﹥绻涢崱妯哄婵炲懐濞€濮婃椽顢�?缂佸鏁婚幃锟犲即閵忥紕鍘繝鐢靛仜閻忔繃淇婇悾�?€妫い鎾跺Т娴滈箖鏌曢崶褍顏い銏℃礋閿燂拷?闁靛繈鍩勯崬铏圭磽閸屾瑦绁板鏉戞憸閺侇噣骞掗弴鐘辫埅闂備浇宕垫慨鏉懨洪妶鍛傜喐绻濋崶褏鍔﹀銈嗗笂閻掞箑鐣风仦鐐弿濠电姴鍟妵婵撴嫹?閿熻姤娲�?〃濠傤潖閼姐倕顥氶悗锝庝簽閸旂敻姊婚崒娆掑厡?闁诲孩绋堥弲婊呮崲濞戞瑧绡€闁告剬鍛暰闂佽�?�╃粙鎺椻€﹂崶鈺佸К闁�?�屽墴濮婃椽骞栭悙鎻掑闂佸憡鏌ㄩˇ鐢哥嵁韫囨拋娲敂閸涱亝�?�奸梻浣告啞缁嬫垿鏁冮敂鍓х＝婵ǹ鍩栭悡鏇㈠箹濞ｎ剨鎷�??閿熶粙宕ú顏呯厽??闂佸府绲介～蹇曠磼濡顎撻梺鍛婄☉閿曘倝寮抽崼婵冩�?妞ゆ梻銆嬪銉х磽瀹ュ拑韬鐐插暣閹粓鎸婃竟鈹垮姂閺屽秹宕崟鑸垫暰闂佸搫鎷嬫禍顏勵潖濞差亜绠伴幖杈剧悼閻ｉ潧顪冮妶蹇撶槣闁搞劋鍗抽�?�娆掔疀閹绢垱鏂€闂�?潻鎷�??閿熺晫绠�???闂傚倷鑳剁划顖濇懌閻熸粍婢橀崯鎾€�?弮鍫晝闁挎梻鏅崢浠嬫⒑閹稿孩纾甸柛�?�崌閿燂拷???婵☆偅绻堝畷娲倷閸濆嫮顓洪梺鎸庢⒒缁垶寮查埡鍛拺閿燂拷?????闂佺ǹ锕ラ幐鎯р枎閵忋�?�鍋ㄩ柛娑樑堥幏娲⒑閸涘﹦鈽夐柨鏇樺劤娴滃憡�?�肩€涙鍘介梺鍐叉惈閿曘�?�鎮�?敃鍌涚厪闁糕剝娲滈ˇ锕傛煃鐠囨煡鍙勬鐐达耿�?�曟﹢鎳犻崹娑樹壕闁割煈鍠掗弨浠嬫煟閹邦厽缍戦柣蹇ョ畵閺岋綁鎮㈤弶鎴犱紙濡ょ姷鍋涚换妯虹暦椤愶箑�?嬮敓锟�????濠碉紕鍋戦崐鏍ь潖婵犳艾纾婚柟鎹愵嚙閸氬綊鏌嶈閸撴瑩鍩為幋锔藉€烽柤纰卞墯閸曢箖姊虹粙鍖℃敾缂佽鐗嗛悾宄懊洪鍕姦濡炪�?�甯婇梽宥嗙濠婂牊鐓欓悗鐢登规禒锕傛�?�濮橆厽�?嬮柡�?€鍠栧畷娆撳Χ閸℃浼�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁€ｅ☉銏犵妞ゆ牗绋戞禒濂告⒑濮瑰浄鎷�??閿熶粙宕归浣侯洸鐟滅増甯楅悡娆撴煟閹寸倖鎴犱焊閻㈠憡鐓曢柡鍌濇硶閸╋綁鏌熼绛嬫畼闁瑰弶鎸抽敓锟�???闁藉嫬銈稿铏圭矙閸ф寮版繛瀛樼矋閸庣厧螞閻斿娓婚柕鍫濇婢ч亶鏌涚€ｎ偆娲撮柟顕嗘�??閿熻В�?介悗锝庝簽椤�?劕鈹戦悜鍥╃У闁告挻鐟︽穱濠囨嚃閳哄啰锛滈梺缁樏幖顐�?触閸︻厾纾奸弶鍫涘妼濞搭喗銇勯姀锛勬噧闁宠閰ｉ幃娆擃敆閸屾簽銉╂⒒娴ｇ瓔鍤欓悗娑掓櫊閹虫繃銈ｉ崘銊幯呯磼鐎ｎ偒鍎ユ繛鍏肩墬缁绘稑顔忛鑽ゅ嚬闂佹悶鍊栫敮锟犲蓟閺囥垹閱囨繝闈涙搐閺呬粙姊洪幐搴ｇ畵闁诡喖娼￠幃鐑藉箥閸愯尙澧梻渚婃嫹?閿熻棄鑻晶浼存煕閹烘挸绗掗柍璇叉唉缁犳盯寮撮悢鍓插晭濠电姷鏁搁敓锟�??婵炰匠鍥ㄥ亱闁告侗鍘搁弻锔姐亜韫囨挾澧涢柛�?�у墲缁绘盯宕卞Ο鍏煎櫘缂備礁顑呴�?�鐑藉蓟閿濆棙鍎熼柕寰涢铏庢繝娈垮枛閿曘劌鈻嶉敐澶婄疅闁圭虎鍠栫粈瀣亜閹伴潧浜濇い銉ヮ儏閳规垿鎮╅锝咁€忛梺鍛婃礀閻忔岸鎮块敓锟�?閹鈻撻崹顔界亶闂佺粯鎼换婵嬫偘閿燂�??瀵粙濡搁敓锟�?椤庢捇姊洪棃鈺佺槣闁告鍘ч锝夊箮閼恒儮鎷绘繛杈剧秬濞咃絿鏁☉娆戠闁告瑥顦辨晶纰夋嫹?閿熻姤娲�?崝姗€濡甸幇鏉跨闁规儳鐡ㄩ鐔兼⒒娴ｈ姤纭堕柛锝忕畵閿燂拷??????
        .ren(backend_dcache_ren),
        .wen(backend_dcache_wen),
        .writen(backend_dcache_writen),
        .vaddr(backend_dcache_addr),
        .write_data(backend_dcache_write_data),

        //trans_addr to dcache
        .ret_data_paddr(ret_data_paddr),
        .duncache_en(duncache_en),

        .dcacop_en(dcacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),
        .cache_axi_write_pre_ready(cache_axi_write_pre_ready),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹瑩寮堕崹顕呭殭闂傚�?�鍊搁崐鐑芥倿閿曞�?�绠栭柛顐ｆ�?绾惧潡鏌ｉ幋鐑嗙劷妞も晛寮剁换婵囩節閸屾粌顤€闂佺ǹ楠哥粔褰掑蓟閿濆绠ｉ柣鎰�?暞缁秶绮嬪鍛牚闁割偆鍠撻崣鍡涙⒑閸濆嫬鏆欐繛鏉戝€垮畷闈涒枎閹存柨浜炬繛鍫濈仢濞呮﹢鏌涢敐蹇曠М鐎殿喖顭烽崹鎯х暦閸ャ劍鐣烽梺璇插嚱缂嶅棝宕滃☉婧惧徍闂傚倸鍊峰ù鍥敋閺嶎厼绐楅柟鐑橆殔閻ょ偓绻濇繝鍌氭灓闁绘帊绮欓悡顐﹀炊閵娿�?�绻�?梺杞扮閸燁垶濡甸崟顖氱�?闁宠桨鑳舵禒濂告⒒婵犲繒鐣垫慨濠傤煼瀹曟帒顫濋钘変壕闁绘垼濮ら崵鍕煕閹捐尙顦﹂柛銊︾箖閵囧嫰寮介顫捕缂備胶濮抽崡鎶藉蓟閻斿吋鈷掗悗鐢登规俊浠嬫⒑缁嬫鍎忔い鎴濐�?瀵鎮㈤崗纭锋�??閿熻姤銇勯幒鍡椾壕婵犫拃灞界仸闁哄本鐩俊鍫曞幢濡⒈妲归梻浣告惈閺堫剟鎯勯鐐靛祦闁搞儺鍓﹂弫鍥煟濮�?棗鏋涘ù鐙呯畵濮婄粯鎷呯粙娆炬闂佺ǹ顑嗙敮妤冪矉�?�ュ鏁傞柛顐ｇ箚閹芥洖鈹戦悙鏉戠仧闁糕晛�?�板顐�?礃椤旂晫鍘梺鍓插亝缁诲啴宕冲ú顏呯厽闊洤娴风粣鏃€鎱ㄦ繝鍐┿仢鐎规洏鍔嶇换娑㈠箳濠靛懘鍋楅梺璇″枟閿氭い顐ｇ箞椤㈡﹢鎮╅锝嗘殼婵犵數濮烽弫鍛婃叏閺夋嚚娲晝閸屾氨锛欐俊鐐差儏缁ㄥ爼宕戦幘缁樺仭闁哄顑欏Λ宀勬⒑閸濄儱校闁绘濮撮悾宄扳堪閸喎浜遍梺鍓插亝缁海绮诲鑸碘拺闂傚牊绋撴晶鏇熺箾鐏炲偊鎷�??閿熶粙鎮ф惔銊︹拻濞达絿鐡旈崵鍐煕閻樺磭澧电€规洘鍔欓獮鏍ㄦ媴閻熼鎮ｉ梻浣虹帛閸ㄧ厧螞閸曨垽缍栭柛娑樼摠閻撳繘鏌涢锝囩畺闁革�?濮ら敓锟�????閻㈩垱甯￠垾鏃堝礃椤斿槈褔鏌涢埄鍏︽岸骞忔繝姘拺闁告繂瀚刊濂告煕鐎ｎ亷宸ラ柣锝囧厴閿燂拷?闁靛牆鎳庣粣娑欑�?閻㈤潧孝閻庢凹鍣ｉ�?�娆撳即閵忥紕鍘告繝銏ｆ硾閿曪附鏅堕弴鐑嗙唵鐟滃繘寮查銈呭灊闁哄啫鐗滈弫鍡椕归敐鍛�?�缂併劏顕ч�?�鍐Χ閸℃顫囬梺绯曟櫅鐎氼剙宓勯梺褰掓？閻掞箓鎮￠悢鍏肩叆婵犻潧妫欓崳瑙勪繆閹绘帩鐓奸柡宀嬬秮閺佹劙宕卞▎鎴犳澖闁诲氦顫夊ú婊堝窗閺嶎叏鎷�?閿熻棄螖閸涱厾锛滃┑顔斤供閸撴盯顢樻總鍛娾拻閿燂�??????闂佺粯甯粻鎾崇暦閺囥垹�?冮悷浣疯兌閹虫捇锝炲┑鍫熷磯闁惧繒娅㈢槐顕€姊虹拠鎻掑毐缂傚秴妫濆畷鎶筋�??鐎殿噮鍋婂畷鎺楁倷鐎电ǹ骞堟俊鐐€栭崝锕傚磻閸曨剚娅犻柟娈垮枤绾惧ジ鎮楅敐搴濈敖缂佺姳鍗抽弻宥囨喆閸曨偆浼岄梺璇″枓閺呮繄妲愰幒鎳崇喐绻濆顓熸婵犵绱曢崑鎴�?磹閺嶎厼鍨傞柣銏⑶圭粻鐘绘煙闁箑鍘存俊鎻掔墦閺岋綁濮€??闂佺粯甯掗悘姘跺Φ閸曨垰绠抽柟瀛樼箥娴犻箖姊洪幎鑺ユ暠闁搞劌婀卞Σ鎰板箻鐎涙ê顎撴繝娈垮枟閸╁牊绂嶅┑瀣疄闁靛ň鏅涢悙濠冦亜閹哄秷鍏岄柛妯圭矙濡懘顢曢姀鈥愁槱闂佸搫琚崝鎴濈暦椤愶附鍊绘俊顖炴櫜缁ㄥ姊洪棃娑氱畾闁糕晛�?�伴獮�?�偐閸愭彃绨ユ繝鐢靛█濞佳兾涢鐑嗙劷闁冲搫鍊舵禍婊堟煙閹屽�??闂佽�?�╂穱鍝勎涢崟顖氱厴闁硅揪闄勯崐鐑芥煠閹间焦娑ф繛鎳峰懐纾藉ù锝囨嚀缁茬粯绻�?????闁伙絿鍏樺鎾閻樻爠鍐剧唵閻犺櫣灏ㄥ銉╂煙椤栨粌浠辨慨濠冩そ閺屽懘鎮欓懠璺侯伃婵犫拃鍐憼闁�?�究鍔嶇换婵嬪礃閳瑰じ铏庢俊銈囧Х閸嬬偤鎮ч悩璇茬畺婵犲﹤鐗嗛悙濠囨煏婵炲灝鍔撮敓锟�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楃€广儱娲ら崹婵囩箾閸℃ɑ灏紒鐘崇墱閹叉悂寮崼婵堢暫闂佸啿鎼崯顖ゆ�??閿熻姤宀搁弻娑樷枎韫囷絾楔闂�?€炲苯澧婚柛鎾跺枎椤繐煤椤忓懎浠梺鍝勵槸缁ㄩ亶骞愰崘顏嗙＝濞撴艾娲ゅ▍姗€鏌涢妸銊︾【妞ゆ洩缍佸濠氬Ψ閵壯屽晣濠电偠鎻徊钘夛�?�闁�?秴鐭楅柛鈩冪⊕閳锋垹绱撴担鐧告嫹???闂備胶枪閿曘倕锕㈤柆宥呯劦妞ゆ帊鑳堕崯鏌ユ煙???
        .rdata(dcache_rdata),
        .rdata_valid(dcache_backend_rdata_valid),    
        .dcache_ready(dcache_ready),  

    //to write BUS
        .dev_wrdy(dev_wrdy_to_cache),      
        .cpu_wen(dcache_wen),        
        .cpu_waddr(dcache_awaddr),      
        .cpu_wdata(dcache_wdata),      
    //to Read Bus
        .dev_rrdy(dev_rrdy_to_cache),       
        .cpu_ren(dcache_ren),        
        .cpu_raddr(dcache_araddr),      
        .dev_rvalid(dcache_rvalid),     
        .dev_rdata(dcache_axi_data_block),
        .ren_received(dcache_ren_received),
    //duncache to cache_axi
        .uncache_rvalid(duncache_rvalid),
        .uncache_rdata(duncache_rdata),
        .uncache_ren(duncache_ren),
        .uncache_raddr(duncache_raddr),

        .uncache_write_finish(duncache_write_finish),
        .uncache_wen(duncache_wen),
        .uncache_wstrb(duncache_wstrb),
        .uncache_wdata(duncache_wdata),
        .uncache_waddr(duncache_waddr)  
    );
        
    addr_trans u_addr_trans(
        .clk(aclk),
        .rst(rst),
        .data_vaddr(backend_dcache_addr),
        .csr_da(csr_da),
        .csr_pg(csr_pg),
        .csr_dmw0(csr_dmw0),
        .csr_dmw1(csr_dmw1),
        .csr_plv(csr_plv),
        .ret_data_paddr(ret_data_paddr),
        .uncache_en(duncache_en)
    );

    axi_interface u_axi_interface(
        .clk(aclk),
        .rst(rst),
    //connected to cache_axi
        .cache_ce(axi_ce_o),
        .cache_wen(axi_wen),   
        .cache_wsel(axi_wsel),      
        .cache_ren(axi_ren),         
        .cache_raddr(axi_raddr),
        .cache_waddr(axi_waddr),
        .cache_wdata(axi_wdata),
        .cache_rready(axi_rready),    
        .cache_wvalid(axi_wvalid),     
        .cache_wlast(axi_wlast),      
        .wdata_resp_o(axi_wdata_resp),    
    
        .cache_brust_type(cache_brust_type),  
        .cache_brust_size(cache_brust_size),
        .cacher_burst_length(axi_rlen),
        .cachew_burst_length(axi_wlen),

        .arid(arid),       
        .araddr(araddr),      
        .arlen(arlen),      
        .arsize(arsize),
        .arburst(arburst),
        .arlock(arlock),   
        .arcache(arcache),   
        .arprot(arprot),   
        .arvalid(arvalid),       
        .arready(arready),         
    //R闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨圭粻璇裁归敐鍫綈闁靛洦绻冮妵鍕閳╁喚妫冮悗瑙勬磸閸�?垿銆佸Ο琛℃斀闁割偆鍠愬В搴ㄦ⒒閸屾熬鎷�??閿熶粙宕愭搴ｇ�???妤犵偞鐗犻�?�鏇氱秴闁搞儺鍓欑粻銉︺亜閺冨�?�鍤€濞存粌澧界槐鎺懳旀担琛℃濠电偞娼欓崐鍨嚕椤愶絿绡€闁搞儯鍔庨崢鎾绘偡濠婂嫮鐭掔€规洘绮撻幃銏＄附婢跺绋佺紓鍌氬€烽悞锕佹懌婵犳鍨遍幐鎶藉蓟閵堝绠掗柟鐑樺灥婵垽姊洪棃娑欘棞闁挎洦浜滈～蹇撁洪鍜佹闂佸啿鎼崯鎷屽€寸紓鍌氬€烽懗鑸垫叏閻㈢ǹ绠查柛銉墯閸嬫ɑ銇勯弮鍥ㄧ�????婵犵數鍋為崹鍫曟偡閿燂拷?閳诲秹濮€閵堝棌鎷洪柣鐘充航閸斿苯鈻嶉幇鐗堢厵闁告垯鍊栭敓锟�????
        .rid(rid),
        .rdata(rdata),   
        .rresp(rresp),    
        .rlast(rlast),           
        .rvalid(rvalid),       
        .rready(rready),
        .rdata_o(axi_rdata),
        .rdata_valid_o(axi_rdata_valid),         
    //AW闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔閹虫捇鈥�?????妞ゅ繐鎳忓畷鎶芥⒑濞茶骞栨俊顐ｇ箞瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻�???婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；婵炴垟鎳為崶顒佸仺缂佸�?�ч悗顒勬⒑閻熸澘鈷旂紒顕呭灦瀹曟垿骞囬悧鍫㈠幘缂佺偓婢樺畷顒佹櫠缂佹ü绻嗛柤纰卞墮閸樺瓨鎱ㄦ繝鍕笡闁瑰嘲鎳樺畷銊︾節閸愩劌澹嶇紓鍌氬€风粈渚€顢栭崟顓燁偨婵﹩鍓涢弳锕傛煏韫囥儳纾挎い鈺冨厴閹鏁愭惔婵堟晼闂佹寧绋掗惄顖氼潖閾忚宕夐柕濞垮劜閻忎焦绻濆▓鍨灓闁轰礁顭烽獮鍐晸閻樿尙顦ㄥ銈嗘⒒閺咁偊宕㈤崡鐐╂斀闁绘绮☉褎淇婇锝庢疁妞ゃ垺妫冮、鏃堝醇閻斿搫骞堥梻浣瑰缁诲�?�骞婇幇顔剧煋婵炲樊浜濋敓锟�????閻庯綆鍓涢敍鐔兼⒑闁偛鑻晶鍓х磼閸欏銇濈€殿喗褰冮埞鎴﹀醇閵忋垹绠甸梻浣告惈閸燁偊鎮ф繝鍥ㄥ亗婵炴垶鍩冮崑鎾诲礂婢跺﹣澹曢梻渚婃嫹?閿熻棄鑻晶杈炬�??閿熻姤娲戦崡鍐差嚕娴犲鏁囬柣妯垮皺閵堬箓姊绘担渚敯闁规椿浜炵划濠氬箣閻樺�?绗夊┑鐐村灟閸ㄦ椽鍩涢幒妤佺厱妞ゆ劑鍊曢弸鏃堟煃椤栨稒绀冮柕鍥у瀵剟宕归鍛棯缂傚�?�鑳剁划顖滄崲閸曨垰绐楀┑鐘蹭迹閻旇铏圭磼濡偐效闂傚倸鍊烽敓锟�??濡炪倖鍨甸幊姗€鐛繝鍌ゆ建闁�?�屽墮椤曪綁顢曢敓锟�??缁€鍐┿亜閺冨�?�鎷℃繛鐓庯躬濮婃椽妫冨☉姘暫闂佺娅曢幑鍥嵁濡ゅ懎鍗抽柕蹇婃�?�閹锋椽姊洪崨濠勭畵閻庢凹鍙冨畷鎺楀Ω閳哄倻鍘遍梺闈浨归崕宕囩矓濞差亝鐓涢悘鐐电摂閸庢棑鎷�??閿熻姤娲栭悥鍏间繆濮濆矈妲鹃梺浼欑畱閻楁挸顫忔繝姘＜婵ê宕敓锟�?缂傚倷绀�?鍡欐暜閻愰潧鍨濆┑鐘叉搐閻撴盯鏌涚仦鍓ф噮缂佺姵鑹鹃—鍐Χ閸℃顫囬梺绋匡攻濞叉绮嬮幒鎴斿牚闁告洍鏅欑花璇差渻閵堝懐绠伴悗姘煎墴�?�娊鏁愰崨顏呮杸闂佺偨鍎辩壕顓㈠春????闁哄洦锚婵倹銇勯姀锛勨�??闁硅偐琛ラ崜婵嬪汲椤忓牊鈷掗敓锟�??????闂佺厧鍟挎晶搴ㄥ礆閹烘鏁嶉柣鎰綑娴滈亶姊洪崫鍕偍闁搞劎鎳撳ú璺ㄧ磽閸屾瑧顦︽い鎴濇椤㈡牕鈻庨幘鍐叉優闂佸搫娲㈤崹娲磻閿濆鐓曢柕澶涚到婵″潡鏌曢崼婵堟憼濞ｅ洤锕獮鎾诲箳閺傛鏉哥紓鍌欒兌缁垳鎹㈤崘顏呭床婵犻潧顑呯壕鍏兼叏濡厧甯跺┑锛勫厴濮婃椽宕妷銉︾€鹃梺璇�?�枛閸婃悂锝炶箛鏃傜瘈婵﹩鍓涢敍婊冣攽閻愬弶顥為柛鏃€顨婃俊鍫曞级鎼存挻鏂€闂佺粯鍔曞Ο濠偽ｇ憴鍕闁肩⒈鍓欓弸搴ㄦ煟閿濆洤鍘存鐐查叄閹崇偤濡烽敂鐣屽絿闂傚倷鑳舵灙闁哄牜鍓欓～婵嬪Ω閳哄﹥鏅╅梺绯曞墲缁嬫帡鍩涢幋锔藉仯闁诡厽甯掓俊鍏肩箾閸涱喖濮嶉柡宀€鍠栧畷娆撳Χ????
        .awid(awid),     
        .awaddr(awaddr),  
        .awlen(awlen),    
        .awsize(awsize),   
        .awburst(awburst),
        .awlock(awlock),   
        .awcache(awcache),
        .awprot(awprot),   
        .awvalid(awvalid),        
        .awready(awready),        
    //W闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔閹虫捇鈥�?????妞ゅ繐鎳忓畷鎶芥⒑濞茶骞栨俊顐ｇ箞瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻�???婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；婵炴垟鎳為崶顒佸仺缂佸�?�ч悗顒勬⒑閻熸澘鈷旂紒顕呭灦瀹曟垿骞囬悧鍫㈠幘缂佺偓婢樺畷顒佹櫠缂佹ü绻嗛柤纰卞墮閸樺瓨鎱ㄦ繝鍕笡闁瑰嘲鎳樺畷銊︾節閸愩劌澹嶇紓鍌氬€风粈渚€顢栭崟顓燁偨婵﹩鍓涢弳锕傛煏韫囥儳纾挎い鈺冨厴閹鏁愭惔婵堟晼闂佹寧绋掗惄顖氼潖閾忚宕夐柕濞垮劜閻忎焦绻濆▓鍨灓闁轰礁顭烽獮鍐晸閻樿尙顦ㄥ銈嗘⒒閺咁偊宕㈤崡鐐╂斀闁绘绮☉褎淇婇锝庢疁妞ゃ垺妫冮、鏃堝醇閻斿搫骞堥梻浣瑰缁诲�?�骞婇幇顔剧煋婵炲樊浜濋敓锟�????閻庯綆鍓涢敍鐔兼⒑闁偛鑻晶鍓х磼閸欏銇濈€殿喗褰冮埞鎴﹀醇閵忋垹绠甸梻浣告惈閸燁偊鎮ф繝鍥ㄥ亗婵炴垶鍩冮崑鎾诲礂婢跺﹣澹曢梻渚婃嫹?閿熻棄鑻晶杈炬�??閿熻姤娲戦崡鍐差嚕娴犲鏁囬柣妯垮皺閵堬箓姊绘担渚敯闁规椿浜炵划濠氬箣閻樺�?绗夊┑鐐村灟閸ㄦ椽鍩涢幒妤佺厱妞ゆ劑鍊曢弸鏃堟煃椤栨稒绀冮柕鍥у瀵剟宕归鍛棯缂傚�?�鑳剁划顖滄崲閸曨垰绐楀┑鐘蹭迹閻旇铏圭磼濡偐效闂傚倸鍊烽敓锟�??濡炪倖鍨甸幊姗€鐛繝鍌ゆ建闁�?�屽墮椤曪綁顢曢敓锟�??缁€鍐┿亜閺冨�?�鎷℃繛鐓庯躬濮婃椽妫冨☉姘暫闂佺娅曢幑鍥嵁濡ゅ懎鍗抽柕蹇婃�?�閹锋椽姊洪崨濠勭畵閻庢凹鍙冨畷鎺楀Ω閳哄倻鍘遍梺闈浨归崕宕囩矓濞差亝鐓涢悘鐐电摂閸庢棑鎷�??閿熻姤娲栭悥鍏间繆濮濆矈妲鹃梺浼欑畱閻楁挸顫忔繝姘＜婵ê宕敓锟�?缂傚倷绀�?鍡欐暜閻愰潧鍨濆┑鐘叉搐閻撴盯鏌涚仦鍓ф噮缂佺姵鑹鹃—鍐Χ閸℃顫囬梺绋匡攻濞叉绮嬮幒鎴斿牚闁告洍鏅欑花璇差渻閵堝懐绠伴悗姘煎墴�?�娊鏁愰崨顏呮杸闂佺偨鍎辩壕顓㈠春????闁哄洦锚婵倹銇勯姀锛勨�??闁硅偐琛ラ崜婵嬪汲椤忓牊鈷掗敓锟�??????闂佺厧鍟挎晶搴ㄥ礆閹烘鏁嶉柣鎰綑娴滃崬鈹戦悩璇у伐闁绘妫濆畷鎺楀Ω瑜庨崰鎰版煛閸愩劎澧涢柡鍛�?閺岋綁骞囬敓锟�?椤ｆ娊鏌ｉ妶鍌氫壕濠电姷鏁搁崑鐐哄垂閸洘鍋￠柨鏇炲€哥壕鎸庛亜韫囨挾澧涢柣鎾跺枛閺岋綁寮幐搴㈠枑闂佺懓鍟块崯鎾箖閿燂拷?椤繈鎮℃惔鈽嗘骄濠电姰鍨奸～澶娒洪悢纭锋嫹?閿熻棄鈽夐姀鈽呮�??閿熺晫绱掗娆炬綈閻庢艾銈稿濠氬磼閿燂�???閹间焦鍋嬪┑鐘叉处閸ゅ嫰鏌涢埄鍐ㄦ惛濞存粌缍婇弻鐔兼倻濡櫣浠奸梺鎸庣�?�閸犳牕顫忓ú顏勪紶闁告洦鍣鍫曟⒑缁嬪灝顒㈤柣鎿勬�??閿熺晫鏆﹂柟鎵椤ュ牊绻涚壕�?�彧婵☆偄鍟村顐�?箛閺夊灝绐涘銈嗘尵閸犳劙顢欐径鎰拻濞达絿鎳撻敓锟�????闂侇剙绉撮崹鍌炴煕瑜庨�?�鍛存嫅閻斿摜绠鹃柟瀵稿€戝璺虹哗濞寸姴顑嗛悡鏇㈡煃閳轰礁鏋ゆ繛鍫涘灩闇夐柣鎾虫捣閻掑憡鎱ㄦ繝鍛仩缂侇喗鐟╁畷绋课旀繛鎯т壕婵°倕鍟扮壕鑲╃磽娴ｅ顏堟倶閺夋垟�?介柨娑樺閺嗩剨鎷�?閿熻姤娲滈崰鏍€佸☉銏℃櫜闁糕剝蓱閻濇繈姊婚崒娆掑厡缂侇噮鍨甸幗顐︽偡濠婂嫭绶查柛鐔告尦閹即顢欓柨顖氫壕闁挎繂楠搁弸鐔兼煃闁垮鐏╃紒杈ㄦ尰閹峰懏鎱ㄩ幋锝呬汗婵炲棎鍨介弻鍡楊吋閸℃瑥骞堥梻浣虹帛閿氱痪缁㈠弮婵℃挳骞掗弮鍌滐紲濡炪倖姊归娆撳吹濞嗘挻鐓冮柦妯侯樈濡叉悂鎽堕敐澶嬧拺闁割煈鍣崕娑欑箾閸忓吋鈷愮紒缁樼箞閹粙妫冨☉妤冩崟婵犵妲呴崑鍛存偡閳轰胶鏆︽繝闈涱儏閿燂�??濡炪倖鎸鹃崰鎰枍閵忋�?�鈷戦悹鎭掑妼濞呮劙鏌�????
        .wid(wid),     
        .wdata(wdata),  
        .wstrb(wstrb),    
        .wlast(wlast),          
        .wvalid(wvalid),       
        .wready(wready),         
    //闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔閹虫捇鈥�?????妞ゅ繐鎳忓畷鎶芥⒑濞茶骞栨俊顐ｇ箞瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻�???婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；婵炴垟鎳為崶顒佸仺缂佸�?�ч悗顒勬⒑閻熸澘鈷旂紒顕呭灦瀹曟垿骞囬悧鍫㈠幘缂佺偓婢樺畷顒佹櫠缂佹ü绻嗛柤纰卞墮閸樺瓨鎱ㄦ繝鍕笡闁瑰嘲鎳樺畷銊︾節閸愩劌澹嶇紓鍌氬€风粈渚€顢栭崟顓燁偨婵﹩鍓涢弳锕傛煏韫囥儳纾挎い鈺冨厴閹鏁愭惔婵堟晼闂佹寧绋掗惄顖氼潖閾忚宕夐柕濞垮劜閻忎焦绻濆▓鍨灓闁轰礁顭烽獮鍐晸閻樿尙顦ㄥ銈嗘⒒閺咁偊宕㈤崡鐐╂斀闁绘绮☉褎淇婇锝庢疁妞ゃ垺妫冮、鏃堝醇閻斿搫骞堥梻浣瑰缁诲�?�骞婇幇顔剧煋婵炲樊浜濋敓锟�????閻庯綆鍓涢敍鐔兼⒑闁偛鑻晶鍓х磼閸欏銇濈€殿喗褰冮埞鎴﹀醇閵忋垹绠甸梻浣告惈閸燁偊鎮ф繝鍥ㄥ亗婵炴垶鍩冮崑鎾诲礂婢跺﹣澹曢梻渚婃嫹?閿熻棄鑻晶杈炬�??閿熻姤娲戦崡鍐差嚕娴犲鏁囬柣妯垮皺閵堬箓姊绘担渚敯闁规椿浜炵划濠氬箣閻樺�?绗夊┑鐐村灟閸ㄦ椽鍩涢幒妤佺厱妞ゆ劑鍊曢弸鏃堟煃椤栨稒绀冮柕鍥у瀵剟宕归鍛棯缂傚�?�鑳剁划顖滄崲閸曨垰绐楀┑鐘蹭迹閻旇铏圭磼濡偐效闂傚倸鍊烽敓锟�??濡炪倖鍨甸幊姗€鐛繝鍌ゆ建闁�?�屽墮椤曪綁顢曢敓锟�??缁€鍐┿亜閺冨�?�鎷℃繛鐓庯躬濮婃椽妫冨☉姘暫闂佺娅曢幑鍥嵁濡ゅ懎鍗抽柕蹇婃�?�閹锋椽姊洪崨濠勭畵閻庢凹鍙冨畷鎺楀Ω閳哄倻鍘遍梺闈浨归崕宕囩矓濞差亝鐓涢悘鐐电摂閸庢棑鎷�??閿熻姤娲栭悥鍏间繆濮濆矈妲鹃梺浼欑畱閻楁挸顫忔繝姘＜婵ê宕敓锟�?缂傚倷绀�?鍡欐暜閻愰潧鍨濆┑鐘叉搐閻撴盯鏌涚仦鍓ф噮缂佺姵鑹鹃—鍐Χ閸℃顫囬梺绋匡攻濞叉绮嬮幒鎴斿牚闁告洍鏅欑花璇差渻閵堝懐绠伴悗姘煎墴�?�娊鏁愰崨顏呮杸闂佺偨鍎辩壕顓㈠春????闁哄洦锚婵倹銇勯姀锛勨�??闁硅偐琛ラ崜婵嬪汲椤忓牊鈷掗敓锟�??????闂佺厧鍟挎晶搴ㄥ礆閹烘鏁嶉柣鎰綑娴滈亶姊洪崫鍕偍闁搞劎鎳撳ú鍧楁⒒娴ｅ摜绉烘俊顐㈡健閹偤鏁冮崒姘憋紱濠殿喗銇涢崑鎾绘煛鐏炶濮傞柟顔哄€濆畷鎺戔槈????闂備浇顕х€涒晠顢欓弽顓炵獥闁哄洨濮撮崹婵囩箾閸℃ê濮冪紒璇叉閺岀喖姊荤€电ǹ濡介梺鍝勬噺缁捇寮诲☉銏犵闁告劦浜欓搹搴ㄦ⒑闂堟稓澧曟い锔垮嵆閸╂盯骞掗幊銊ョ秺閺佹劙宕奸悤浣峰摋闂佹眹鍩勯崹閬嶆儎椤栫偛钃熸繛鎴欏灩缁秹鏌熼幆褍顣抽柡鍡愬€濋幃妤冩喆閸曨剛顦ㄧ紓渚囧枛閻�?�宕洪姀鈩冨劅闁靛ǹ鍎抽鎾绘⒑閸涘﹤濮€闁哄懏绮岄埢宥夊幢濞戞瑢鎷绘繛杈剧秬婵倗娑甸崼鏇熺厱闁挎繂绻掗悾鍨殽閻愯尙绠婚柡浣规崌閿燂拷???
        .bid(bid),      
        .bresp(bresp),    
        .bvalid(bvalid),        
        .bready(bready)         
    );

    cache_AXI u_cache_AXI(
        .clk(aclk),
        .rst(rst),    // low active

    //icache read
        .inst_ren_i(icache_ren),
        .inst_araddr_i(icache_araddr),
        .inst_rvalid_o(icache_rvalid),
        .inst_rdata_o(icache_rdata),
        .icache_ren_received(icache_ren_received),
        .icache_flush_flag_valid(icache_flush_flag_valid),

    //dcache read
        .data_ren_i(dcache_ren),
        .data_araddr_i(dcache_araddr),
        .data_rvalid_o(dcache_rvalid),
        .data_rdata_o(dcache_axi_data_block),
        .dcache_ren_received(dcache_ren_received),

    //dcache write
        .data_wen_i(dcache_wen),
        .data_wdata_i(dcache_wdata),
        .data_awaddr_i(dcache_awaddr),
        .data_bvalid_o(dcache_bvalid),

        .cache_axi_write_pre_ready(cache_axi_write_pre_ready),

    //ready to cache
        .dev_rrdy_o(dev_rrdy_to_cache),
        .dev_wrdy_o(dev_wrdy_to_cache),

    //uncache to dcache
        .duncache_ren_i(duncache_ren),
        .duncache_raddr_i(duncache_raddr),
        .duncache_rvalid_o(duncache_rvalid),
        .duncache_rdata_o(duncache_rdata),

        .duncache_wen_i(duncache_wen),
        .duncache_wstrb(duncache_wstrb),
        .duncache_wdata_i(duncache_wdata),
        .duncache_waddr_i(duncache_waddr),
        .duncache_write_resp(duncache_write_finish),

    //AXI communicate
        .axi_ce_o(axi_ce_o),
        .axi_wsel_o(axi_wsel),   // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ら敓锟�?闁秴鐒垫い鎺戝€归敓锟�??闁诲孩鍑归崣鍐ㄧ暦�?�曞洤顥氶悗锝冨妺濮规姊洪崷顓炲妺闁搞劌缍婂畷鎰版倷閻戞ê浠┑鐘诧工閿燂拷???闁诲孩顔栭崰妤呭箖閸屾凹鍤曞ù鐘差儛閺佸洭鏌ｉ弬鎸庢儓妤犵偞鍔欏缁樻媴鐟欏嫬浠╅梺绋垮瘨閸ㄨ泛鐣烽弴銏＄劶閿燂拷?????闂備礁鍟块幖顐﹀疮閹殿喖顥氬┑鍌氭啞閻撴瑩姊�????鐎殿喚鍋撶换娑㈠醇閻旇櫣鐓夐敓锟�??????闁伙絾绻堥敓锟�?妞ゆ帒�?�粣妤呮煛瀹ュ骸骞栫紒鐘崇墱閹叉悂寮捄銊︽婵犻潧鍊搁幉锟犲磻閸曨垱鐓曟繝闈涙椤忊晜绻涢崼娑樺姦婵﹤顭峰畷鎺戔枎閹搭厽袦闂備胶顢婇婊呮崲濠靛棛鏆﹂柛锔诲幗閸犲棝鏌�????鐎殿喖娼″娲捶椤撯剝顎楅梺鍝ュУ閻楃娀骞冮垾鎰佹建闁�?�屽墴�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戠紒瀣儥閸庢劙鏌涢敓锟�??閻熲晠鐛�?崘銊庢棃宕ㄩ鐔风ザ婵＄偑鍊栭幐楣冨磹椤愶箑顫呴幒铏濠婂牊鐓忓鑸电☉椤╊剛绱掗悩鎰佺劷缂佽鲸甯�?蹇涘Ω閿燂拷?闂夊秹姊洪悷鏉挎Щ闁硅櫕锚閻ｇ兘顢曢敓锟�?缁€瀣棯閻�?煫顏呯????闁�?�屽墴�?�曠喖顢楅崒姘疄闂傚�?�绶氶敓锟�??闂佺ǹ瀛╂繛濠傜暦濞差亝鏅查柛銉到娴滅偓绻涢崼婵堜虎闁哄绋掗妵鍕敇閻樻彃骞嬮悗娈垮櫘閸嬪﹪鐛�?崶顒夋晣闁绘劗鏁搁悰顔尖攽閻樺灚鏆╁┑顔碱嚟?濮樺崬鍘寸€规洏鍎靛畷顭掓嫹?閿熻姤菤閹风粯绻涙潏鍓ф偧闁硅櫕鎹囬�?�姘堪閸涱垳锛滈柣鐘叉处瑜板啴鍩€閿燂�??濞硷繝鎮伴钘夌窞濠电偟鍋撻～宥夋⒑闂堟稓绠冲┑顔惧厴椤㈡瑩骞掗弮鍌滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋為崰姗堟�??閿熻姤娲忛崹浠嬬嵁閺嶃劍濯撮柛蹇擃槹鐎氬ジ姊绘担鍛婂暈缂佸鍨块弫鍐晲閸ヮ煈鍋ㄩ梻渚囧墮缁夌敻鎮￠弴銏＄厽婵☆垵顕ф晶顖涚箾閸喓鐭岄柍褜鍓濋～澶娒洪敓锟�?瀹曟繂鈻庨幘璺虹ウ闂佹悶鍎洪崜姘跺磻鐎ｎ喗鐓曟い鎰Т閻忊晜顨ラ悙鏉戝婵﹨娅ｉ幑鍕Ω閵夛妇褰氶梻浣烘嚀閿燂�?????闂傚倷娴囬褔宕欓悾�?€绀婇柛鈩冪☉缁€鍫熺箾閹存瑥鐏柛搴★躬閺屾盯顢曢悩鎻掑闂佺ǹ锕﹂弫濠氬箖瀹勬壋鏋庨煫鍥ㄦ惄娴犲墽绱撴担鎻掍壕闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄被鍔岄埞鎴�?醇濠靛懐鎹曟俊銈嗩殢娴滄瑩宕￠崘鑼殾闁绘挸绨堕弨浠嬫�?�閿濆簼绨奸柡鍡�?邯濮婂宕掑▎鎺戝帯缂備緡鍣�?崹璺侯嚕婵犳艾惟闁崇懓绨遍崑鎾诲礃閳哄�?�鍔呴梺闈涒康闂勫嫬鈻嶉�?銈嗏拺閻犳亽鍔屽▍鎰版煙????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌￠敓锟�??閸犳牠骞冭瀹曞ジ鎮㈤崫鍕闂傚�?�绀�?幉锟犲垂鐟欏嫭鍙忛柟缁㈠枛閻撴﹢鏌熸潏楣冩�?�闁稿鍔欓幃妤呭捶椤撶倫銏°亜閵夛妇绠樼紒杈ㄦ尰閹峰懘宕�?????闂備焦鎮堕崝�?勬偉閻撳寒鍤曞┑鐘宠壘鎯熼梺鍐叉惈閸婂憡绂嶉悙鐑樷拺缂佸�?�у﹢鎵磼鐎ｎ偄鐏存い銏℃閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧櫢鎷�??閿熻棄�?�崳纾嬨亹閹烘垹鍊為悷婊冾�?瀵悂寮介鐔哄幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柟閭�?弾濞堟粓鏌�?�畝瀣瘈鐎规洖鐖奸崺鈩冩媴閹绘帊澹曢梺鎸庣箓閹冲危閸儲鐓忛煫鍥ㄦ礀鍟稿銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛鈩兠弳妤佺節濞堝灝鏋ら柛蹇斍瑰Λ鐔奉渻閵堝棛澧紒瀣尵�?�囧焵椤掑嫭鈷戞慨鐟版搐閻忓弶绻涙担鍐插暟閹姐儱鈹戦悩鍨毄闁稿鐩幆鍥ㄥ閺夋垹锛欏┑鐘绘涧椤戝懐绮婚鐐寸厵閺夊牓绠栧顕€鏌涚€ｎ亜顏柡灞剧缁犳稑顫濋鎸庣潖闂備礁鎲￠敃鈺傜濠靛牊宕叉繝闈涱儐閸嬨劑姊婚崼鐔衡棩闁瑰鍏樺铏圭矙濞嗘儳鍓遍梺鐟版啞閹�?�宕洪姀鐙€鍚嬪璺猴工閼板灝鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶愭涧闇夋繝濠傚閻帗銇勯姀鈩冾棃妞ゃ垺锕㈤敓锟�??闁挎稑�?�獮鎰版⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掔€ｎ亞鍙€婵犮垼鍩栭崝鏍偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺撳暈闁靛洤�?�伴、鏇㈡晲閸モ晝鍘滈柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟�??楠炪垽鏌嶉崫鍕舵�??閿熺晫绮婇鐣岀瘈闁汇垽娼у暩闂佽桨鐒﹂幃鍌氱暦閹存績妲堥柕蹇婃櫆閺咁亜顪冮妶鍡樺蔼闁搞劌缍婂畷鎺�?Ω瑜庨崰鎰節闂堟侗鍎忕紒鐙€鍨堕弻銊╂偆閸屾稑顏�??闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧闁绘柨妫欓幈銊ヮ渻鐠囪弓澹曢梻浣瑰缁诲嫰宕戦悩鐢典笉婵炴垯鍨瑰Λ姗€鎮归崶顏勭处闁哥姴锕娲嚒閵堝懏鐎洪梻鍌氬缁夌懓鐣烽幇鏉跨闁归潧鐏曢崗鐐�?�曘劑顢欑憴鍕伖闂傚�?�绶氬浼欐�??閿熻棄鐭傚畷銏＄附缁嬭法顦柣搴秵閸撴稓澹曟總鍛婂仯闁搞儯鍔岀徊濠氭煛閸☆厾绉�?柟绋匡躬閹垽宕楅懖鈺佸箰闁诲骸绠嶉崕杈殽閹间胶宓佹俊銈呮噺閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵娿儳顑傞梺閫炲苯澧剧紓宥呮瀹曘垽鎮剧仦鎯у幑闂佸憡鎸烽懗鍓佸婵傚憡鐓熸俊顖濇閿涘秹鏌涘▎灞戒壕闂傚�?�绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌℃径�?�闁绘柨鍚嬮幆鐐烘⒑椤愶絿鈯曢柛瀣噹閳规垿鏁嶉崟顐℃澀闂佺ǹ锕ラ悧鏇犲弲闂佸啿鎼崯鎵矆婵犲偊鎷�?閿熻棄顫濋敐鍛闂備線娼уΛ鏃傛濮橆剦鍤曢柟缁㈠枛椤懘鏌嶉埡浣告殲闁绘繃鐗犻敓锟�???闁�?�屽墰閸嬫盯鎳熼娑欐珷闁规鍠氱壕鍏笺亜閺傚灝鈷旈悽顖涚�?�缁辨帞绱掑Ο鑲╃暤濡炪�?�鍋呯换鍫ャ€侀敓锟�??閹晠骞撻幒鏃傛澖闂傚�?�鍊搁崐宄懊归崶顒婄稏濠㈣泛锕﹂弳锔戒繆椤栫偞锛熼柣鎺戯攻缁绘盯宕卞Ο璇差伇闂佹悶鍎洪崜姘跺疾濠婂牊鐓曢煫鍥ㄦ�?鐢埖銇�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楅柡鍥╁枑閸欏繘鏌曢崼婵囧仾濡わ箒娉曢敓锟�??濠电偞鍨堕�?�鍥晬閻斿吋鈷掑�?�姘搐婢ь喚绱掓径妯烘珝??濡炪倖甯婇悞锕偹�?????闁哄洨鍣﹂懓鎸庛亜閵忥紕鎳囩€规洖寮剁粩鐔碱敍濮橆厼顦╅梺缁樻尰濞茬喖寮诲澶婄厸濞达絿枪缁犺顪冮妶鍛闁绘妫楁晥闁告瑥顦换鍡涙煏閸繂顏柛蹇撶灱缁辨帡鍩�??闁稿鎸荤换婵嬫偨闂堟稐绮堕梺缁橆殔濡繈骞冨Ο琛℃斀閿燂�??????閿燂�?????缂佸鏁婚幃锟犲即閻旇櫣顔曢梺绯曞墲椤ㄥ牏绮绘导瀛樼厸闁糕剝顭囬幊鍕煏閸パ冾伃鐎殿喗鎸抽�?�鏃堝幢濞呯儤绮撻幃妤冩喆閸曨剛顦ㄩ梺鎸庡哺濡焦寰勯幇顓ㄦ�??閿熶粙鏌ㄥ┑鍡欏嚬缂併劏妫勯…鑳檨闁搞劏娉涢～蹇曠磼濡顎撶紓浣割儐椤戞瑥螞瀹€鍕拺缂佸顑欓崕蹇斾繆椤愶絿绠撻柣锝夋敱鐎靛ジ寮堕幋鐙€鍟嬮梺鑽ゅТ濞诧箒銇愰崘顔肩；鐎广儱顦伴埛鎴︽煕閹剧懓鐨洪柛妯荤洴閺屾冻鎷�??????闂佺懓绠嶉崹钘夌暦閸楃偐妲堟繛鍡樺灥楠炴姊绘担鍝ョШ闁稿锕畷婊冾潩鐠鸿櫣鍘洪梺鍝勬储閸ㄦ椽鎮￠弴銏犵閺夊牆澧界壕璺ㄧ磼閻樺樊鐓奸柡�?€鍠栭�?�娆戠驳鐎ｎ偆鏉�????闁哄洨鍋熺粔鐑樸亜閵忊剝�?嬮敓锟�??闂傚嫬娲敓锟�???婵﹦绮幏鍛驳鐎ｎ亝鐣伴梻浣告憸婵敻骞戦崶褏鏆︾憸鐗堝笚鐎电姴顭跨捄鐑樻拱婵炲牓绠栧娲箰鎼达絺妲堥柣搴㈠嚬閸犳碍绂嶉幖浣瑰仺闁汇垻鏁搁敍婊堟⒑闂堟胆褰掑磿椤栫偛鐒垫い鎺戯攻閿燂拷?

    //AXI read
        .rdata_i(axi_rdata),
        .rdata_valid_i(axi_rdata_valid),
        .axi_ren_o(axi_ren),
        .axi_rready_o(axi_rready),
        .axi_raddr_o(axi_raddr),
        .axi_rlen_o(axi_rlen),

    //AXI write
        .wdata_resp_i(axi_wdata_resp),  // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔閹虫捇鈥�?????妞ゅ繐鎳忓畷鎶芥⒑濞茶骞栨俊顐ｇ箞瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻�???婵犲痉甯嫹?閿熻姤鎱ㄩ悜钘夌；婵炴垟鎳為崶顒佸仺缂佸�?�ч悗顒勬⒑閻熸澘鈷旂紒顕呭灦瀹曟垿骞囬悧鍫㈠幘缂佺偓婢樺畷顒佹櫠缂佹ü绻嗛柤纰卞墮閸樺瓨鎱ㄦ繝鍕笡闁瑰嘲鎳樺畷銊︾節閸愩劌澹嶇紓鍌氬€风粈渚€顢栭崟顓燁偨婵﹩鍓涢弳锕傛煏韫囥儳纾挎い鈺冨厴閹鏁愭惔婵堟晼闂佹寧绋掗惄顖氼潖閾忚宕夐柕濞垮劜閻忎焦绻濆▓鍨灓闁轰礁顭烽獮鍐晸閻樿尙顦ㄥ銈嗘⒒閺咁偊宕㈤崡鐐╂斀闁绘绮☉褎淇婇锝庢疁妞ゃ垺妫冮、鏃堝醇閻斿搫骞堥梻浣瑰缁诲�?�骞婇幇顔剧煋婵炲樊浜濋敓锟�????閻庯綆鍓涢敍鐔兼⒑闁偛鑻晶鍓х磼閸欏銇濈€殿喗褰冮埞鎴﹀醇閵忋垹绠甸梻浣告惈閸燁偊鎮ф繝鍥ㄥ亗婵炴垶鍩冮崑鎾诲礂婢跺﹣澹曢梻渚婃嫹?閿熻棄鑻晶杈炬�??閿熻姤娲戦崡鍐差嚕娴犲鏁囬柣妯垮皺閵堬箓姊绘担渚敯闁规椿浜炵划濠氬箣閻樺�?绗夊┑鐐村灟閸ㄦ椽鍩涢幒妤佺厱妞ゆ劑鍊曢弸鏃堟煃椤栨稒绀冮柕鍥у瀵剟宕归鍛棯缂傚�?�鑳剁划顖滄崲閸曨垰绐楀┑鐘蹭迹閻旇铏圭磼濡偐效闂傚倸鍊烽敓锟�??濡炪倖鍨甸幊姗€鐛繝鍌ゆ建闁�?�屽墮椤曪綁顢曢敓锟�??缁€鍐┿亜閺冨�?�鎷℃繛鐓庯躬濮婃椽妫冨☉姘暫闂佺娅曢幑鍥嵁濡ゅ懎鍗抽柕蹇婃�?�閹锋椽姊洪崨濠勭畵閻庢凹鍙冨畷鎺楀Ω閳哄倻鍘遍梺闈浨归崕宕囩矓濞差亝鐓涢悘鐐电摂閸庢棑鎷�??閿熻姤娲栭悥鍏间繆濮濆矈妲鹃梺浼欑畱閻楁挸顫忔繝姘＜婵ê宕敓锟�?缂傚倷绀�?鍡欐暜閻愰潧鍨濆┑鐘叉搐閻撴盯鏌涚仦鍓ф噮缂佺姵鑹鹃—鍐Χ閸℃顫囬梺绋匡攻濞叉绮嬮幒鎴斿牚闁告洍鏅欑花璇差渻閵堝懐绠伴悗姘煎墴�?�娊鏁愰崨顏呮杸闂佺偨鍎辩壕顓㈠春????闁哄洦锚婵倹銇勯姀锛勨�??闁硅偐琛ラ崜婵嬪汲椤忓牊鈷掗敓锟�??????闂佺厧鍟挎晶搴ㄥ礆閹烘鏁嶉柣鎰綑娴滈亶姊洪崫鍕偍闁搞劎鎳撳ú鍧楁⒒娴ｅ摜绉烘俊顐㈡健閹偤鏁冮崒姘憋紱濠殿喗銇涢崑鎾绘煛鐏炶濮傞柟顔哄€濆畷鎺戔槈????闂備浇顕х€涒晠顢欓弽顓炵獥闁哄洨濮撮崹婵囩箾閸℃ɑ灏柍褜鍏涚欢姘嚕閹绢喖顫呴柍銉ュ帠缁ㄥ姊绘担鍝勪壕闁煎綊绠栧畷鎰板箹閿燂拷?婢跺⿴娼╂い鎾跺Х閻﹀牓姊哄Ч鍥х伈婵炰匠鍕浄闁挎洖鍊归悡鏇㈡煏婵炲灝鍔ら柛鈺嬬稻閵囧嫰濮€閳╁啠鎷归柣搴ㄦ涧閵堢ǹ顕ｉ崼鏇炵�???闁告艾鎳忕换娑欐綇閸撗冨煂缂備礁顦靛褔顢氶妷鈺佺妞ゆ牗姘ㄩ敓锟�?婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓熷顐ャ亹閹烘挴鎷绘繛鎾村焹閸嬫挻绻涙担鍐叉瘽閵娾晛鐒�??闁宠鍨块崹楣冩惞椤愩垺鐏庨柣搴ゎ潐濞插繘宕归挊澶屾殾闁靛⿵濡囬敓锟�??闂佸憡娲﹂崣搴ㄥ疮鎼淬劍鈷戦柛婵嗗濡叉悂鏌ｉ敓锟�?濡瑩寮查崼鏇熷�???闁活厽鎸婚妵鍕箳�?�ュ顎栨繛瀛樼矋缁秹濡甸崟顖氱疀闁宠桨鑳堕崝鏉戔攽閳ュ啿绾ч柟顔煎€垮濠氭晲婢跺娅滈梺鍛婁緱閸樻垝绨洪梻鍌欐缁鳖喚寰婇崜褎宕查柛顐ｇ箘閺嗭箓鏌ｉ弮鍌楁嫛闁轰礁妫濋弻娑氫沪閹规劕顥濈紓浣哄О閸庨潧顫忔繝姘＜婵炲棙鍨垫俊浠嬫⒑缁嬪潡顎楅柛鐔锋健濠€浣糕攽椤旇鐟扳枖濞戞艾顥氱憸鐗堝笚閸婄敻鏌ㄥ┑鍡涱€楁繛鍛�?�閺屸剝鎷�????闂佸搫鏈惄顖炪€侀弴銏╂晝闁靛繒濯鍓х磽閸屾瑧顦︽い鎴濇噽閹广垽骞囬弶璺ㄥ幋闂佺鎻梽鍕磻閹邦喚纾藉ù锝堝亗閹达附鐓ユい鎾跺剱濞撳鏌曢崼婵囶棞闁诲繈鍎甸弻鐔兼惞椤愩垹顫岄梺瀹犳椤︾敻骞冮悾宀€鐭欓悹鎭掑妼婵附淇婇悙顏庢嫹?閿熺晫鏁�?敓锟�???濮樼厧寮�?柛鈺傜洴楠炲鎮╅悽纰夌闯濠电偠鎻徊浠嬶綖閺嶎収鏁傞柛娑卞枛�?�潡姊洪幖鐐插姶闁告挻�?搁幃锟犳偄閼测晛褰勯梺鎼炲劘閸斿秹鎮￠妷鈺傜厱婵犻潧鐗嗛崝�?�煏閸パ冾�???闂佹剚鍘搁弲婊堝垂瑜版帒绠查柕蹇曞Л閺€浠嬫煕閿燂�??閺呮粓宕撻棃娑辨富闁靛牆妫欑亸鎵磼鐎ｎ偄绗ч柍褜鍓氭穱鍝勎涢崟顖氱厴闁硅揪闄勯崐鐑芥煠閹间焦娑ф繛鎳峰懐纾藉ù锝囨嚀缁茬粯绻�?????闁伙絿鍏樺鎾閻樻爠鍐剧唵閻犺櫣灏ㄥ銉╂煙椤栨粌浠辨慨濠冩そ閺屽懘鎮欓懠璺侯伃婵犫拃鍐憼闁�?�究鍔嶇换婵嬪礃閳瑰じ铏庢俊銈囧Х閸嬬偤鎮ч悩璇茬畺婵犲﹤鐗嗛悙濠囨煏婵炲灝鍔撮敓锟�????闂傚倸鍊峰ù鍥р枖閺囥垹绐楃€广儱娲ら崹婵囩箾閸℃ɑ灏紒鐘崇墱閹叉悂寮崼婵堢暫闂佸啿鎼崯顖ゆ�??閿熻姤宀搁弻娑樷枎韫囷絾楔闂�?€炲苯澧婚柛鎾跺枎椤繐煤椤忓懎浠梺鍝勵槸缁ㄩ亶骞愰崘顏嗙＝濞撴艾娲ゅ▍姗€鏌涢妸銊︾【妞ゆ洩缍佸濠氬Ψ閵壯屽晣濠电偠鎻徊钘夛�?�闁�?秴鐭楅柛鈩冪⊕閳锋垹绱撴担鐧告嫹???闂備胶枪閿曘倕锕㈤柆宥呯劦妞ゆ帊鑳堕崯鏌ユ煙???
        .axi_wen_o(axi_wen),
        .axi_waddr_o(axi_waddr),
        .axi_wdata_o(axi_wdata),
        .axi_wvalid_o(axi_wvalid),
        .axi_wlast_o(axi_wlast),
        .axi_wlen_o(axi_wlen)
    );


    wire [101:0] data1;
    wire [101:0] data2;
    wire valid1;
    wire valid2;
    wire [101:0] debug_data_out;
    wire debug_valid_out;

    assign data1 = {debug_wb_we1,debug_reg_addr1,debug_wdata1,debug_inst1,debug_pc1};
    assign data2 = {debug_wb_we2,debug_reg_addr2,debug_wdata2,debug_inst2,debug_pc2};
    assign valid1 = debug_wb_valid1;
    assign valid2 = debug_wb_valid2;
/*
    debug_FIFO debug
    (
        .clk(aclk),
        .rst(rst),
        .valid1(valid1),
        .data1(data1),
        .valid2(valid2),
        .data2(data2),
        .data_out(debug_data_out),
        .valid_out(debug_valid_out)
    );
*/
    assign debug0_wb_pc = 0;  
    assign debug0_wb_rf_wen = 0;
    assign debug0_wb_rf_wnum = 0;
    assign debug0_wb_rf_wdata = 0;

endmodule