`timescale 1ns / 1ps
`include "defines.vh"

module core_top(
    input  wire        aclk,
    input  wire        aresetn,
    input  wire [ 7:0] intrpt, 
    //AXI interface 
    //read reqest
    output wire [ 3:0] arid,
    output wire [31:0] araddr,
    output wire [ 7:0] arlen,
    output wire [ 2:0] arsize,
    output wire [ 1:0] arburst,
    output wire [ 1:0] arlock,
    output wire [ 3:0] arcache,
    output wire [ 2:0] arprot,
    output wire        arvalid,
    input  wire        arready,
    //read back
    input  wire [ 3:0] rid,
    input  wire [31:0] rdata,
    input  wire [ 1:0] rresp,
    input  wire        rlast,
    input  wire        rvalid,
    output wire        rready,
    //write request
    output wire [ 3:0] awid,
    output wire [31:0] awaddr,
    output wire [ 7:0] awlen,
    output wire [ 2:0] awsize,
    output wire [ 1:0] awburst,
    output wire [ 1:0] awlock,
    output wire [ 3:0] awcache,
    output wire [ 2:0] awprot,
    output wire        awvalid,
    input  wire        awready,
    //write data
    output wire [ 3:0] wid,
    output wire [31:0] wdata,
    output wire [ 3:0] wstrb,
    output wire        wlast,
    output wire        wvalid,
    input  wire        wready,
    //write back
    input  wire [ 3:0] bid,
    input  wire [ 1:0] bresp,
    input  wire        bvalid,
    output wire        bready,

    // debug
    
    input           break_point,    //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剟鎮块敓锟???閺岋絽螖閳ь剟鎮ц箛鏇犱笉濡わ絽鍟悡鍐喐濠婂牆绀堟慨妯块哺�?�曞弶绻涢幋娆忕仼缂佺姴顭烽弻娑㈠箛椤掍讲鏋欓梺鍝勬閸ㄨ棄顫忓ú顏呯劵闁绘劘灏�??锟戒即鏌ㄩ悤鍌涘�????闂傚倷绶￠崜娆戠矓鐎电ǹ顥氬┑鐘崇閻撶喖鏌￠崘銊︽悙濞存粌婀遍埀顒冾潐閹搁娆㈠璺鸿摕婵炴垯鍨瑰敮濡炪倖姊婚崢褔锝為敓�??????濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柣鏂垮悑閻撴盯鏌涢幇鈺佸缂佷讲鏅犻弻娑㈠Χ閸℃瑦鍣伴梺鍝勬湰缁嬫垼鐏掔紓鍌欑劍閿氶柛鐐差�?濮婃椽宕崟顕呮蕉闂佸憡鏌ㄩ惌鍌炲春閵夛箑绶炲┑鐐灮閸犳劗绮悢纰辨晬婵炴垵宕弫宕囩磽閸屾熬�????閿熶粙宕愭搴㈩偨闁跨喓濮寸粣妤呮煛瀹ュ骸骞楅柣鎾亾闂備焦瀵х换鍌炈囬崡鐐垫殼濞撴埃鍋撻柡锟??鍠栭獮鎴�?箛闂堟稒顔勭紓鍌欒兌婵數绮欓幒�???桅闁告洦鍠氶敓锟???闂佸湱鍋撻幆灞轿涢妷褏纾藉ù锝堟鐢盯鏌涢妸銉т虎妞ゎ偄绻�?幖鍦喆閸曨偅鐎梻浣告啞濞诧附绂嶉敐澶婃槬闁告稑鐡ㄩ埛鎴犵磼鐎ｎ偄顕滈柛鐐差槺缁辨帡顢氶埀顒傜不閺嶃劋绻嗛柣銏⑶圭粻娑欍亜閹达絽袚妞ゎ偄绉瑰娲濞戞氨顔婃繝娈垮枤閸忔﹢濡撮敓�????瀹曨煉锟???閿熻姤菤閹锋椽姊洪崨濠勨槈闁挎洏鍊栭幈銊╁醇閵忥�??锟芥瀾闂佸搫顦悘婵嬪汲閻斿吋鐓欙拷?锟藉嫰鍋婇崕鏃撴�??閿熺瓔鍠栭�?�閿嬩繆閻戣姤鏅滈柟顖嗗啯杈堟繝鐢靛Х閺佹悂宕戦悙鍝勫瀭闁割偅娲嶉�?顒婄畵�?�曞爼顢楁担绯曞亾閸噮娓婚悗锝庝簼閹癸絿鐥崜褍甯堕摶鐐烘煟閿燂拷?閻楀繒绮婚幘鍨涘亾濞堝灝娅橀柛锝忕秮瀵鍩勯崘鈺侊�??锟介柣鐔哥懃鐎氼剛澹曢幎鑺モ拺閺夌偞澹嗛崝宥夋煙閻熺増鍠橈拷?锟筋噮鍋婇獮妯肩磼濡粯�??????1闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛顐ｆ礀绾惧鏌曟繛鐐珔缁炬儳娼￠弻锛勪沪鐠囨彃濮曢梺绋款儐閿曘垽寮婚敓锟?????0
    input           infor_flag,     //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剟鎮块敓锟???閺岋絽螖閳ь剟鎮ц箛鏇犱笉濡わ絽鍟悡鍐喐濠婂牆绀堟慨妯块哺�?�曞弶绻涢幋娆忕仼缂佺姴顭烽弻娑㈠箛椤掍讲鏋欓梺鍝勬閸ㄨ棄顫忓ú顏呯劵闁绘劘灏�??锟戒即鏌ㄩ悤鍌涘�????闂傚倷绶￠崜娆戠矓鐎电ǹ顥氬┑鐘崇閻撶喖鏌￠崘銊︽悙濞存粌婀遍埀顒冾潐閹搁娆㈠璺鸿摕婵炴垯鍨瑰敮濡炪倖姊婚崢褔锝為敓�??????濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柣鏂垮悑閻撴盯鏌涢幇鈺佸缂佷讲鏅犻弻娑㈠Χ閸℃瑦鍣伴梺鍝勬湰缁嬫垼鐏掔紓鍌欑劍閿氶柛鐐差�?濮婃椽宕崟顕呮蕉闂佸憡鏌ㄩ惌鍌炲春閵夛箑绶炲┑鐐灮閸犳劗绮悢纰辨晬婵炴垵宕弫宕囩磽閸屾熬�????閿熶粙宕愭搴㈩偨闁跨喓濮寸粣妤呮煛瀹ュ骸骞楅柣鎾亾闂備焦瀵х换鍌炈囬崡鐐垫殼濞撴埃鍋撻柡锟??鍠栭獮鎴�?箛闂堟稒顔勭紓鍌欒兌婵數绮欓幒�???桅闁告洦鍠氶敓锟???闂佸湱鍋撻幆灞轿涢妷褏纾藉ù锝堟鐢盯鏌涢妸銉т虎妞ゎ偄绻�?幖鍦喆閸曨偅鐎梻浣告啞濞诧附绂嶉敐澶婃槬闁告稑鐡ㄩ埛鎴犵磼鐎ｎ偄顕滈柛鐐差槺缁辨帡顢氶埀顒傜不閺嶃劋绻嗛柣銏⑶圭粻娑欍亜閹达絽袚妞ゎ偄绉瑰娲濞戞氨顔婃繝娈垮枤閸忔﹢濡撮敓�????瀹曨煉锟???閿熻姤菤閹锋椽姊洪崨濠勨槈闁挎洏鍊栭幈銊╁醇閵忥�??锟芥瀾闂佸搫顦悘婵嬪汲閻斿吋鐓欙拷?锟藉嫰鍋婇崕鏃撴�??閿熺瓔鍠栭�?�閿嬩繆閻戣姤鏅滈柟顖嗗啯杈堟繝鐢靛Х閺佹悂宕戦悙鍝勫瀭闁割偅娲嶉�?顒婄畵�?�曞爼顢楁担绯曞亾閸噮娓婚悗锝庝簼閹癸絿鐥崜褍甯堕摶鐐烘煟閿燂拷?閻楀繒绮婚幘鍨涘亾濞堝灝娅橀柛锝忕秮瀵鍩勯崘鈺侊�??锟介柣鐔哥懃鐎氼剛澹曢幎鑺モ拺閺夌偞澹嗛崝宥夋煙閻熺増鍠橈拷?锟筋噮鍋婇獮妯肩磼濡粯�??????1闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛顐ｆ礀绾惧鏌曟繛鐐珔缁炬儳娼￠弻锛勪沪鐠囨彃濮曢梺绋款儐閿曘垽寮婚敓锟?????0
    input  [ 4:0]   reg_num,        //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剟鎮块敓锟???閺岋絽螖閳ь剟鎮ц箛鏇犱笉濡わ絽鍟悡鍐喐濠婂牆绀堟慨妯块哺�?�曞弶绻涢幋娆忕仼缂佺姴顭烽弻娑㈠箛椤掍讲鏋欓梺鍝勬閸ㄨ棄顫忓ú顏呯劵闁绘劘灏�??锟戒即鏌ㄩ悤鍌涘�????闂傚倷绶￠崜娆戠矓鐎电ǹ顥氬┑鐘崇閻撶喖鏌￠崘銊︽悙濞存粌婀遍埀顒冾潐閹搁娆㈠璺鸿摕婵炴垯鍨瑰敮濡炪倖姊婚崢褔锝為敓�??????濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柣鏂垮悑閻撴盯鏌涢幇鈺佸缂佷讲鏅犻弻娑㈠Χ閸℃瑦鍣伴梺鍝勬湰缁嬫垼鐏掔紓鍌欑劍閿氶柛鐐差�?濮婃椽宕崟顕呮蕉闂佸憡鏌ㄩ惌鍌炲春閵夛箑绶炲┑鐐灮閸犳劗绮悢纰辨晬婵炴垵宕弫宕囩磽閸屾熬�????閿熶粙宕愭搴㈩偨闁跨喓濮寸粣妤呮煛瀹ュ骸骞楅柣鎾亾闂備焦瀵х换鍌炈囬崡鐐垫殼濞撴埃鍋撻柡锟??鍠栭獮鎴�?箛闂堟稒顔勭紓鍌欒兌婵數绮欓幒�???桅闁告洦鍠氶敓锟???闂佸湱鍋撻幆灞轿涢妷褏纾藉ù锝堟鐢盯鏌涢妸銉т虎妞ゎ偄绻�?幖鍦喆閸曨偅鐎梻浣告啞濞诧附绂嶉敐澶婃槬闁告稑鐡ㄩ埛鎴犵磼鐎ｎ偄顕滈柛鐐差槺缁辨帡顢氶埀顒傜不閺嶃劋绻嗛柣銏⑶圭粻娑欍亜閹达絽袚妞ゎ偄绉瑰娲濞戞氨顔婃繝娈垮枤閸忔﹢濡撮敓�????瀹曨煉锟???閿熻姤菤閹锋椽姊洪崨濠勨槈闁挎洏鍊栭幈銊╁醇閵忥�??锟芥瀾闂佸搫顦悘婵嬪汲閻斿吋鐓欙拷?锟藉嫰鍋婇崕鏃撴�??閿熺瓔鍠栭�?�閿嬩繆閻戣姤鏅滈柟顖嗗啯杈堟繝鐢靛Х閺佹悂宕戦悙鍝勫瀭闁割偅娲嶉�?顒婄畵�?�曞爼顢楁担绯曞亾閸噮娓婚悗锝庝簼閹癸絿鐥崜褍甯堕摶鐐烘煟閿燂拷?閻楀繒绮婚幘鍨涘亾濞堝灝娅橀柛锝忕秮瀵鍩勯崘鈺侊�??锟介柣鐔哥懃鐎氼剛澹曢幎鑺モ拺閺夌偞澹嗛崝宥夋煙閻熺増鍠橈拷?锟筋噮鍋婇獮妯肩磼濡粯�??????5闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛顐ｆ礀绾惧鏌曟繛鐐珔缁炬儳娼￠弻锛勪沪鐠囨彃濮曢梺绋款儐閿曘垽寮婚敓锟?????0
    output          ws_valid,       //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剟鎮块敓锟???閺岋絽螖閳ь剟鎮ц箛鏇犱笉濡わ絽鍟悡鍐喐濠婂牆绀堟慨妯块哺�?�曞弶绻涢幋娆忕仼缂佺姴顭烽弻娑㈠箛椤掍讲鏋欓梺鍝勬閸ㄨ棄顫忓ú顏呯劵闁绘劘灏�??锟戒即鏌ㄩ悤鍌涘�????闂傚倷绶￠崜娆戠矓鐎电ǹ顥氬┑鐘崇閻撶喖鏌￠崘銊︽悙濞存粌婀遍埀顒冾潐閹搁娆㈠璺鸿摕婵炴垯鍨瑰敮濡炪倖姊婚崢褔锝為敓�??????濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柣鏂垮悑閻撴盯鏌涢幇鈺佸缂佷讲鏅犻弻娑㈠Χ閸℃瑦鍣伴梺鍝勬湰缁嬫垼鐏掔紓鍌欑劍閿氶柛鐐差�?濮婃椽宕崟顕呮蕉闂佸憡鏌ㄩ惌鍌炲春閵夛箑绶炲┑鐐灮閸犳劗绮悢纰辨晬婵炴垵宕弫宕囩磽閸屾熬�????閿熶粙宕愭搴㈩偨闁跨喓濮寸粣妤呮煛瀹ュ骸骞楅柣鎾亾闂備焦瀵х换鍌炈囬崡鐐垫殼濞撴埃鍋撻柡锟??鍠栭獮鎴�?箛闂堟稒顔勭紓鍌欒兌婵數绮欓幒�???桅闁告洦鍠氶敓锟???闂佸湱鍋撻幆灞轿涢妷褏纾藉ù锝堟鐢盯鏌涢妸銉т虎妞ゎ偄绻�?幖鍦喆閸曨偅鐎梻浣告啞濞诧附绂嶉敐澶婃槬闁告稑鐡ㄩ埛鎴犵磼鐎ｎ偄顕滈柛鐐差槺缁辨帡顢氶埀顒傜不閺嶃劋绻嗛柣銏⑶圭粻娑欍亜閹达絽袚妞ゎ偄绉瑰娲濞戞氨顔婃繝娈垮枤閸忔﹢濡撮敓�????瀹曨煉锟???閿熻姤菤閹锋椽姊洪崨濠勨槈闁挎洏鍊栭幈銊╁醇閵忥�??锟芥瀾闂佸搫顦悘婵嬪汲閻斿吋鐓欙拷?锟藉嫰鍋婇崕鏃堟煥閻曞�?�锟?????
    output [31:0]   rf_rdata,       //闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剟鎮块敓锟???閺岋絽螖閳ь剟鎮ц箛鏇犱笉濡わ絽鍟悡鍐喐濠婂牆绀堟慨妯块哺�?�曞弶绻涢幋娆忕仼缂佺姴顭烽弻娑㈠箛椤掍讲鏋欓梺鍝勬閸ㄨ棄顫忓ú顏呯劵闁绘劘灏�??锟戒即鏌ㄩ悤鍌涘�????闂傚倷绶￠崜娆戠矓鐎电ǹ顥氬┑鐘崇閻撶喖鏌￠崘銊︽悙濞存粌婀遍埀顒冾潐閹搁娆㈠璺鸿摕婵炴垯鍨瑰敮濡炪倖姊婚崢褔锝為敓�??????濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柣鏂垮悑閻撴盯鏌涢幇鈺佸缂佷讲鏅犻弻娑㈠Χ閸℃瑦鍣伴梺鍝勬湰缁嬫垼鐏掔紓鍌欑劍閿氶柛鐐差�?濮婃椽宕崟顕呮蕉闂佸憡鏌ㄩ惌鍌炲春閵夛箑绶炲┑鐐灮閸犳劗绮悢纰辨晬婵炴垵宕弫宕囩磽閸屾熬�????閿熶粙宕愭搴㈩偨闁跨喓濮寸粣妤呮煛瀹ュ骸骞楅柣鎾亾闂備焦瀵х换鍌炈囬崡鐐垫殼濞撴埃鍋撻柡锟??鍠栭獮鎴�?箛闂堟稒顔勭紓鍌欒兌婵數绮欓幒�???桅闁告洦鍠氶敓锟???闂佸湱鍋撻幆灞轿涢妷褏纾藉ù锝堟鐢盯鏌涢妸銉т虎妞ゎ偄绻�?幖鍦喆閸曨偅鐎梻浣告啞濞诧附绂嶉敐澶婃槬闁告稑鐡ㄩ埛鎴犵磼鐎ｎ偄顕滈柛鐐差槺缁辨帡顢氶埀顒傜不閺嶃劋绻嗛柣銏⑶圭粻娑欍亜閹达絽袚妞ゎ偄绉瑰娲濞戞氨顔婃繝娈垮枤閸忔﹢濡撮敓�????瀹曨煉锟???閿熻姤菤閹锋椽姊洪崨濠勨槈闁挎洏鍊栭幈銊╁醇閵忥�??锟芥瀾闂佸搫顦悘婵嬪汲閻斿吋鐓欙拷?锟藉嫰鍋婇崕鏃堟煥閻曞�?�锟?????

    output [31:0] debug0_wb_pc,
    output [ 3:0] debug0_wb_rf_wen,
    output [ 4:0] debug0_wb_rf_wnum,
    output [31:0] debug0_wb_rf_wdata

    `ifdef DIFF
    ,
    // difftest
    output [31:0] debug1_wb_pc,
    output [ 3:0] debug1_wb_rf_wen,
    output [ 4:0] debug1_wb_rf_wnum,
    output [31:0] debug1_wb_rf_wdata,
    output [31:0] debug1_wb_inst
    `endif

);

        `ifdef DIFF
    // difftest
    reg             cmt0_valid        ;
    reg             cmt0_cnt_inst     ;
    reg     [63:0]  cmt0_timer_64     ;
    reg     [ 7:0]  cmt0_inst_ld_en   ;
    reg     [31:0]  cmt0_ld_paddr     ;
    reg     [31:0]  cmt0_ld_vaddr     ;
    reg     [ 7:0]  cmt0_inst_st_en   ;
    reg     [31:0]  cmt0_st_paddr     ;
    reg     [31:0]  cmt0_st_vaddr     ;
    reg     [31:0]  cmt0_st_data      ;
    reg             cmt0_csr_rstat_en ;
    reg     [31:0]  cmt0_csr_data     ;

    reg             cmt1_valid        ;
    reg             cmt1_cnt_inst     ;
    reg     [63:0]  cmt1_timer_64     ;
    reg     [ 7:0]  cmt1_inst_ld_en   ;
    reg     [31:0]  cmt1_ld_paddr     ;
    reg     [31:0]  cmt1_ld_vaddr     ;
    reg     [ 7:0]  cmt1_inst_st_en   ;
    reg     [31:0]  cmt1_st_paddr     ;
    reg     [31:0]  cmt1_st_vaddr     ;
    reg     [31:0]  cmt1_st_data      ;
    reg             cmt1_csr_rstat_en ;
    reg     [31:0]  cmt1_csr_data     ;
 
    reg     [ 3:0]  cmt0_wen          ;
    reg     [ 7:0]  cmt0_wdest        ;
    reg     [31:0]  cmt0_wdata        ;
    reg     [31:0]  cmt0_pc           ;
    reg     [31:0]  cmt0_inst         ;
    reg             cmt0_excp_flush   ;
    reg             cmt0_ertn         ;
    reg     [5:0]   cmt0_csr_ecode    ;
    reg             cmt0_tlbfill_en   ;

    reg     [ 3:0]  cmt1_wen          ;
    reg     [ 7:0]  cmt1_wdest        ;
    reg     [31:0]  cmt1_wdata        ;
    reg     [31:0]  cmt1_pc           ;
    reg     [31:0]  cmt1_inst         ;
    reg             cmt1_excp_flush   ;
    reg             cmt1_ertn         ;
    reg     [5:0]   cmt1_csr_ecode    ;
    reg             cmt1_tlbfill_en   ;
    reg     [4:0]   cmt_rand_index    ;

    // to difftest debug
    reg             trap                  ;
    reg     [ 7:0]  trap_code             ;
    reg     [63:0]  cycleCnt              ;
    reg     [63:0]  instrCnt              ;
 
    // from regfile 
    reg     [31:0]  regs_diff[31:0]       ;
    wire    [31:0]  regs_diff_out[31:0]   ;

    // from ctrl
    wire    [`DIFF_WIDTH-1:0] diff0           ;
    wire    [`DIFF_WIDTH-1:0] diff1           ;
    wire    [63:0]  cnt                   ;
  
    // from csr  
    wire    [31:0]  csr_crmd_diff_0       ;
    wire    [31:0]  csr_prmd_diff_0       ;
    wire    [31:0]  csr_ectl_diff_0       ;
    wire    [31:0]  csr_estat_diff_0      ;
    wire    [31:0]  csr_era_diff_0        ;
    wire    [31:0]  csr_badv_diff_0       ;
    wire	[31:0]  csr_eentry_diff_0     ;
    wire 	[31:0]  csr_tlbidx_diff_0     ;
    wire 	[31:0]  csr_tlbehi_diff_0     ;
    wire 	[31:0]  csr_tlbelo0_diff_0    ;
    wire 	[31:0]  csr_tlbelo1_diff_0    ;
    wire 	[31:0]  csr_asid_diff_0       ;
    wire 	[31:0]  csr_save0_diff_0      ;
    wire 	[31:0]  csr_save1_diff_0      ;
    wire 	[31:0]  csr_save2_diff_0      ;
    wire 	[31:0]  csr_save3_diff_0      ;
    wire 	[31:0]  csr_tid_diff_0        ;
    wire 	[31:0]  csr_tcfg_diff_0       ;
    wire 	[31:0]  csr_tval_diff_0       ;
    wire 	[31:0]  csr_ticlr_diff_0      ;
    wire 	[31:0]  csr_llbctl_diff_0     ;
    wire 	[31:0]  csr_tlbrentry_diff_0  ;
    wire 	[31:0]  csr_dmw0_diff_0       ;
    wire 	[31:0]  csr_dmw1_diff_0       ;
    wire 	[31:0]  csr_pgdl_diff_0       ;
    wire 	[31:0]  csr_pgdh_diff_0       ;
    `endif 



    wire rst;
    assign rst = !aresetn;

    wire icache_ren;
    wire [31:0] icache_araddr;
    wire icache_rvalid;
    wire [255:0] icache_rdata;
    wire dcache_ren;
    wire [31:0] dcache_araddr;
    wire dcache_rvalid;
    wire [31:0] dcache_rdata;
    wire [3:0] dcache_wen;
    wire [255:0] dcache_wdata;
    wire [31:0] dcache_awaddr;
    wire dcache_bvalid;

    //AXI communicate
    wire axi_ce_o;
    wire [3:0] axi_wsel;   
    //AXI read
    wire [31:0] axi_rdata;
    wire axi_rdata_valid;
    wire axi_ren;
    wire axi_rready;
    wire [31:0] axi_raddr;
    wire [7:0] axi_rlen;
    wire [255:0] dcache_axi_data_block;

    //AXI write
    wire axi_wdata_resp;
    wire axi_wen;
    wire [31:0] axi_waddr;
    wire [31:0] axi_wdata;
    wire axi_wvalid;
    wire axi_wlast;
    wire [7:0] axi_wlen;
    wire [1:0] cache_brust_type;
    assign cache_brust_type = 2'b01;   
    wire [2:0] cache_brust_size;
    assign cache_brust_size = 3'b010;

    //icache  闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????缂傚倸鍊烽懗鑸垫叏閻㈢ǹ鍨傞柛褎顨呴弰銉╂煏韫囧�????閿熶粙宕￠幎鑺ョ厪闊洢鍎崇壕鍧楁煕濞嗗繑顥㈡慨濠呮缁辨帒螣閼姐�?�妲梺璺ㄥ櫐閿燂拷????????濠电姷鏁告慨鐑斤�??锟介鐐潟闁哄洢鍨圭壕濠氭煙鏉堝墽鐣辩痪鎯х秺閺岋拷?锟筋吋鎼达拷?锟界凹闂佸搫妫欑划鎾诲蓟閻斿吋鍊绘慨�???妫欓悾鍓佺磼閻愵剙鍔ら敓�????闁秴绠熼柟闂寸劍閸嬪鏌涢锝囩畼闁荤喐鐓″娲传閸曨剙娅ら梺璇″枛閸婂灝顕ｆ繝姘╅柍鍝勶�??锟芥禍鐐烘⒑缁嬫寧婀扮紒瀣灴閺佹捇鏁撻敓锟?????闂傚倸鍊搁崐鎼佸磹閹间礁纾癸�??锟藉嫭鍣磋ぐ鎺戠倞妞ゆ帒顦伴弲顏堟偡濠婂啰绠婚柛鈹惧亾濡炪�?�甯婇懗鍫曞煝閹剧粯鐓涢柛娑卞灠瀛濋梺浼欑到閸㈡煡鍩㈡惔銊ョ閻庯絺鏅滈惈蹇涙⒒娴ｅ憡璐￠柛搴涳�??锟藉畷褰掓偨缁嬭法锛涢悗骞垮劚濡稓寮ч埀顒勬煥閻曞�?�锟???????缂傚倷鑳堕搹搴ㄥ储婵傚憡鍋夊┑鍌溓归敓锟????濠碉紕鍋戦崐鏍暜閹烘鏅濋柨鏇烇拷?锟介敓锟???????闂備礁鎼ú銊╁磻閻旇櫣鐭撻柣鎴炃滄禍婊堟煏韫囧ň鍋撻崘鍙夋嚈闁诲氦顫夊ú蹇涘礉閹达讣�????閿熻棄鈻庨幘鏉戞異闂佸啿鎼崯顐λ囬埡鍛拻闁稿本鑹鹃�?顒佹倐�?�曟劖顦版惔銏╁仺濠殿喗枪濞夋盯鎮為崹顐犱簻闁圭儤鍨甸埀�???鎲＄粋鎺戔堪閸喓鍘惧┑鐐跺蔼椤曆囨倶閿熺姵鐓涢柛娑卞幘閸╋綇锟???閿熺瓔鍠栭�?�閿嬩繆閻戣姤鏅滈柟顖嗗啰顔戞繝纰夌磿閸嬫垿宕愰弽顓炵闁割偅娲栭崹鍌氣攽閻樺磭顣查柛�?�ф櫊閺岋綁骞嬮悙鍡樺灴�?�曪�?绠涢幘顖涙杸闂佺粯蓱瑜板啴寮抽悙鐑樼厪闁搞儯鍔庨敓锟????闁荤喐鐟ワ拷?锟筋厾澹曢幖浣圭厱闁哄�?�娉曡�?�闂佺懓绠嶉崹褰掑煘閹寸姭鍋撻敐搴濈敖妞わ缚鍗冲娲濞戞帒鎮嶉柣搴ㄦ涧閼活垶鈥﹂崶锟??绫嶉柛顐ゅ暱閹峰姊虹粙鎸庢拱闁荤啙鍥佸洭鏁傛慨鎰盎闂佽宕樼亸娆撴儗濞嗘垟鍋撳▓鍨灈闁绘牜鍘ч悾鐤亹閹烘繃鏅梺鍛婁緱閸犳氨绮旈悽鍛娾拻闁稿本鑹鹃�?顒傚厴閹虫宕滄担鐟板幑闂佸壊鍋呭ú鏍偪閻愵剛锟??濠电姴鍊绘晶娑㈡煕鎼达拷?锟筋劉闁靛洤瀚板浠嬵敃椤厽鍩涢柣搴ゎ潐閹搁娆㈠璺虹畺婵°�?�鎳忛弲鏌ュ箹缁懓澧查柣蹇撶Ч濮婃椽宕崟锟??娅ょ紓渚囧枟閹瑰洤顕ｆ繝姘櫢闁跨噦�????闁句紮绲介妴鎺戭潩閻撳海浠柛鐔告�?�濮婄粯鎷呴崨濠傛殘闂佺粯顨嗛�?�濠囧箖瑜旈幃鈺侇啅椤旂晫绋佺紓鍌氾�??锟介悞锕佹懌婵犳鍨伴顓犳閹烘垟妲堟慨锟??妫楅崜鏉库攽閻愯尙澧涢柛�???鐟ラ～蹇撁洪鍕獩婵犵數濮村ù鐑藉礉閻戣姤鈷戦柛婵嗗婵ジ鏌涳�??锟筋亷宸ユい鏇秮椤㈡洟鏁傜紒妯绘珨闂備緤锟???閿熻棄鑻晶鎾煟濞戝崬娅嶆鐐村浮閺佹捇鏁撻敓�?????缂備胶濮撮�?�鐑藉蓟閵堝洤鏋堥柛妤冨仜椤偊姊烘导娆戠ɑ闁稿孩濞婇崺鐐哄箣閿旇棄浜圭紓鍌欑劍钃遍梺娆惧弮濮婅櫣绮欓崠鈩冩暰闂佽鍠栭崐鍧楁偘椤旇棄绶為柟閭�?幗濞呫垽姊虹紒妯忣亪宕幐搴ｎ洸婵°�?�鍋撻柍瑙勫灴閹瑩寮堕幋鐘辨埛闂備焦鎮堕崝宥咁渻閽樺鏆﹂柟鎵閸嬨劑鏌涘☉姗堝姛闁告瑥妫楅埞鎴︽偐缂佹ɑ閿┑鈽嗗亝缁诲牓銆�?幘缁樻櫢闁跨噦锟???闂傚洤顦扮换婵囩�?閸屾凹锟??闂佹椿鍘界敮锟犲蓟閳ュ磭鏆嗛悗锝庡墰琚ｇ紓鍌欒兌婵敻鎯勯姘煎殨妞ゆ洍鍋撻柛鈹惧亾濡炪倖甯掗崐鐑芥倿婵犲洦鐓ラ柡鍥╁仜閳ь剙缍婇幃鈥斥槈閵忊槄锟???閿熶粙鏌ｉ幇顔芥毄闁靛棗锕弻娑虫嫹?閿熺瓔鍋呯亸顓㈡煟閿濆洤鍘达�??锟芥洖鐖兼俊鎼佹晜閻愵剚顔曢梻鍌氾拷?锟藉ù鍥敋瑜斿畷娆撴偩閿燂拷?�???濠囨煕閳╁啰鈽夐敓锟???閸喓绠鹃柟瀛樼懃閻忣亪鏌￠崪浣稿⒋闁哄矉缍佸顒勫垂椤�?枻锟???閿熶粙姊洪幎鑺ユ暠闁搞劌鐏濋～蹇撁洪宥嗘櫇闂侀潧鐗嗛幊宥囧垝閸洘鈷戦柛蹇撳悑閵囩喖鏌涢妸�???鎲撅�??锟筋喗鐓″畷濂稿即閻愭妲堕柣鐔哥矊缁绘帗绔熼敓�????????闂備線娼чˇ顓㈠磿閺屻儱闂柣鎴炃滄禍婊堟煏婢诡垰鍟╅幋椋庣磽娴ｄ粙鍝洪悽顖ゆ嫹?閿熺晫鏆﹂柟鐑樺焾濞尖晜鎱ㄩ敐鍡欐嚂闁瑰嚖锟????闁荤喐鐟ワ拷?锟筋厾绮堥埀顒勬⒑闂堟稓澧㈤弸顏呫亜閺囶亞绉鐐达耿椤㈡瑩鎸婃径澶�?泿闂傚�?�鑳堕崑鎾绘嚌妤ｅ啫纾瑰┑鐘宠壘濮瑰弶淇婇妶鍛櫤闁抽攱甯￠弻娑氫沪閸撗勫櫙闂佺ǹ绻愰惌鍌氼嚕閹间緡鏁傞柛鈩冪懅閿涙粎绱撻崒娆戝妽闁挎碍绻涢幖顓炴珝闁哄本鐩崺锟犲磼濠婂嫬鍨遍柣搴ゎ潐濞叉粓宕㈣閸╃偤骞嬮敓锟???�???鍐煃閸濆嫬鏆曠紒銊ョ摠缁绘繈鎮介棃娑楃捕濡炪�?�娲﹂崢浠嬪箞閵娾晛绠绘い鏇炴噺閺呯偤姊虹化鏇炲⒉缂佸甯�?�畷鎴﹀磼閻愬鍘介梺鍝勶拷?锟介悘婵嬪箖閹达附鐓熼柟鎯ь嚟閹冲洦鎱ㄦ繝鍐┿仢妞ゃ垺锕㈡俊姝岊槾闁哄棛锟??濮婅櫣鎷犻懠顒傤唺闂佽法鍣﹂敓锟????闂備礁鎼惌澶岀礊娴ｏ拷?锟界箚闁归棿�?佹儫闂佹寧妫�?濠囧传濡ゅ啰纾介柛灞剧懄缁佹澘顪冮弶鎴炴喐闁轰緡鍣ｉ弫鎾绘偐閼碱剛鏆梻浣哥枃濡椼劎娆㈤敓鐘茬柈闁告侗鍠撴禍婊堟煥閻曞倹锟???闂佺ǹ瀛╂繛濠囩嵁閸愵喖绠ｉ柨鏃囆掗幏缁樼箾鏉堝墽鍒伴柟璇х�?楠炲棝宕奸妷锔惧幗濡炪�?�鎸鹃崕鎰ｉ悜妯圭箚闁告瑥顦慨宥忔嫹?閿熺瓔鍠楅幐鎶藉箖閵忥紕鐟规い鏍ㄧ�?�閵堫偊姊婚崒娆戝妽閻庣瑳鍐炬綎濠电姵鑹鹃敓�????????婵犳鍠楁灙闁糕晜鐗犻幃鈥斥枎閹寸姷锛濇繛杈剧到椤牠顢旈崨顖楁敵濡炪�?�鐗滈崑鐐烘偂閻旂厧绠归弶鍫濆⒔閸掍即鏌涘Ο铏规憼闁�?�究鍔嶇换婵嬪礋椤撶偟顐肩紓鍌欑劍椤ㄥ牓宕伴弽顓熸櫢闁跨噦锟???闂佽法鍣﹂敓�????????濠碉紕鍋戦崐鏍暜閹烘纾归柛娑橈功椤╅攱绻濇繝鍌滃�?闁绘挾濮电换娑㈡嚑妫版繂娈梺璇查獜缁绘繈寮婚敓鐘插窛妞ゆ挾濮撮悡鐔兼�?�鐟欏嫭�?冪紒顔肩箻钘濋悗闈涙憸濡垶鏌熼鍡曠娴狀噣姊洪崫鍕潶闁稿﹥绻堥獮濠傗攽鐎ｎ亞楠囬柣鐘充航閸斿瞼鏁幐搴濈箚闁绘劦浜滈埀顒佸灴�?�曟洟鏌嗗畵銉ユ喘閹晫绮欑捄顭戝晥闂備礁澹婇崑鍛洪敓�????瀹曟劙鎮滈懞銉у幗闂佺懓顕崕鎰版倿娴犲鐓曟俊顖滅帛閸婃劖鎱ㄦ繝鍐┿仢鐎规洏鍔嶇换婵嬪磼濮樺吋缍嗛梻鍌欑閹诧繝寮婚妸鈺傛櫢闁跨噦锟?????濠碉紕鍋戦崐鏍ь啅婵犳艾纾婚柟鎯у绾炬枻锟???閿熷鍎遍幏鎴︾叕椤掑嫭鐓忛柛鈩冩礈缁愭棑锟???閿熺瓔鍠楅幐铏叏閳ь剟鏌嶉妷銊︾彧闁汇�?�鎳樺缁樼瑹閳ь剙顭囪閺佹捇鏁撻敓�?????缂傚倷鑳舵慨鐢稿垂閻㈠壊鏁嬮柨婵嗩槸閸ㄥ倹銇勯弮鍥舵綈闁哄�?�鍋撻梻鍌欑閻ゅ洤螞閸曨�?�娑樜旈崨顕嗘嫹?閿熶粙鏌ㄩ悢鍝勑ｉ柛濠勬暩缁辨帒螖娴ｈ�??妲堥梺鐟板暱缁绘ê鐣烽敓锟???楗即宕楅悙顒侇棃闁轰焦鍔欏畷銊╊敇閻斿壊鍞归梻鍌欒兌缁垶骞愰崼鏇炲�?�濞寸姴顑呴拑鐔哥箾閹存瑥鐏╃紒鐘崇洴閺屾稖绠涢幘�?�樺枑闂佺儵鏅涢柊锝咁潖濞差亜浼犻柛鏇㈡涧閸撻亶姊洪悜鈺傛珦闁搞劏娉涢锝嗙�?濮橆厽娅栭梺鍛婃处娴滄繈宕熼崘顔解拺缂備焦锚婵箓鏌涢幘瀵告创閽樻繈鏌曟繛褍鎳愰敍婵囩箾鏉堝墽绉繛鍜冪悼閺侇喖鈽夐�?锛勫幗闂佸啿鎼敃銈夋�?�閿旂瓔娈介柣鎰絻閺嗘瑩鏌嶇拠鏌ュ弰妤犵偞鐟╁畷锟??鍩￠崒娑氬綅濠电姷鏁搁崑鐘诲箵椤忓棗绶ゅù鐘差儏缁犺銇勯幇鈺嬫嫹?閿熺晫娆㈤妶鍛傛棃鏁愰崨顓熸闂佹娊�?辩敮锟犲蓟濞戞矮娌柛鎾�?嫬娅欓梻浣呵圭换鎰版儗閸屾凹鍤曢柟闂寸贰閺佸倿鏌涘☉鍗炰簵缂併劌顭峰娲偡閹殿喗鎲肩紓浣筋嚙閸熸潙鐣烽搹顐ゎ浄閻庯綆鍋嗛崢鎾绘偡濠婂嫮鐭掞�??锟芥洘绮岄～婵嬫嚋闂堟稑�?????闁诲氦顫夊ú鈺冩崲濠靛棛鏆︽俊顖欒閸熷懏銇勯弬鍨�?�妞ゆ挸娼�?�娲嚒閵堝憛銏＄箾鐠囇冾洭缂侇喖锕鍫曞箠缁涘湱绉拷?锟芥洖銈搁幃銏ゅ礈娴ｈ櫣鏆板┑锛勫亼閸婃牠鎮у⿰鍫濈；闁绘劕鎼弸�???寮堕崼娑樺Ω濞存粍绮嶉妵鍕箛閳轰胶浼勯悗娑欑箞濮婄尨�????閿熺晫濯鎰版煕閵娿儲鍋ラ柕鍡曠閳诲酣骞嬮悩鐑╂敽闂佽鍑界紞鍡涘磻閸℃稑姹查柕澶嗘櫆閳锋帒霉閿濆牊顏犻悽顖涚⊕閵囧嫰濡搁妷�???娅ｉ柧鑽ゅ仦缁绘盯宕卞Ο璇茬缂備胶濮烽崑銈夊蓟閺囩喓绠鹃柛顭戝枛婵鈹戦埄鍐ㄧ祷闁绘锕﹂幑銏犫槈閵忕姴鑰垮┑鈽嗗灥濞咃絾绂掗悡搴富闁靛牆妫欓埛鎰箾閼碱剙鏋涳�??锟筋喖顭烽弫鎰板幢濡搫濡抽梻浣瑰缁诲倸螞濞嗗警鎺�?礋椤栨稓鍘搁柣搴到閿燂�??闂侇収鍨堕弻鐔碱敊閼姐�?�鐓撳銈冨灪缁嬫垿锝炲┑�?�闁绘劙娼ч獮妤呮⒒閸屾瑦绁版い鏇熺墵瀹曟澘螖閸涱�?鍋撻崘顔煎窛閺夊牆澧界粙蹇撯攽閻樼粯娑фい鎴炲姍�?�偊宕堕浣哄幗闂佸搫鍊癸�??锟窖囧箚閸儲鐓曢柕鍫濇缁楁艾菐閸パ嶈含闁诡噯�???????闂傚倷鑳舵灙妞ゆ垵鎳愰埀顒佸嚬閸ｏ綁鐛幋锟??顫呴柕鍫濇噽閿燂�??婵＄偑鍊栧濠氬储瑜旈幃鍧楀箚瑜夐弨浠嬫煥濞戞ê顏╁ù婊愭嫹???缂傚倸鍊烽懗鍓佸垝椤栫偛�?夋俊銈呮噹閻掑灚銇勯幒宥囶槮闁搞値鍓熼弻娑樜熼幁鎺戜划闂佽鍣ｇ粻鏍涢崘銊㈡闁告鍋為崐顖炴⒒娴ｅ憡鍟炵紒顔肩墦閹偤鏁傞崗鐓庮�??闂佽法鍠曞Λ鍕儗閸屾凹娼栨繛宸簼椤ュ牊绻涢幋鐐跺妞わ絽鎼埞鎴﹀煡閸℃ぞ绨奸梺鑽ゅ暀閸曨収娲搁梺褰掓？閻掞箓宕戦妸鈺傜厱婵炴垶锕崝鐔兼煕閿燂拷?娴滃爼寮婚敐鍡樺劅妞ゆ牗绮庢牎闂備胶枪椤戝懎螞濡ゅ啫寮查梻浣告贡閾忓酣宕板Δ鍛亗闁绘柨鎽滅粻楣冩煙鐎涙绠撻柤绋跨秺閺屸槄锟???閿熷鍔岄埀顒佺箞�?�顓奸崼顐ｏ�??锟介梻浣告啞閹稿爼宕濇惔锝嗩潟闁绘劕鎼獮銏＄箾閹寸儐鐒介柣娑栧劚閳规垶骞婇柛濠冩礋楠炲﹥鎯旈妸�???浜楅梺鍝勬储閸ㄦ椽鎮″▎鎾崇骇闁割偁鍎抽悾鐑樹繆缂併垹娅嶉柡灞剧〒閳ь剨缍嗛崜娆愮墡缂傚�?�鑳剁划顖炴儎椤栫偟宓侀悗锝庡枟閺呮煡鏌涢埄鍐噧婵炴嚪鍥ㄢ拺閻犲洦褰冮銏ゆ煟閺冩垵澧存鐑囨�???闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖鎮ч崼鐔哄嚒闂佹悶鍔岄崐鍦崲濠靛顥堟繛鎴炵懃缁愭盯姊虹紒妯肩畵闁绘牕銈稿濠氭晸閻樿尙鍊為梺闈涱槶閸庤櫕绂掓ィ鍐┾拺闁规儼濮ら弫閬嶆偨椤栥�?�锟??鐎殿喛顕ч埥澶婎潩椤愶絽濯伴梻浣告啞閹稿棝宕熼锝囧蒋闂傚倷娴囧畷鍨叏閻㈢ǹ绀夐柟鐑橆殔閿燂拷?闂佽鍎煎Λ鍕嫅閻斿摜绠鹃柟瀛樼懃閻忊晝绱掗悩宸吋闁诡喗顨婂Λ鍐ㄢ槈濞嗗繑娈�?梻锟??娼荤紞鍡涘窗濮樿鲸顫曢柟鎯ь嚟閻熷綊鏌涢妷鎴濆娴滆埖绻濈喊妯活潑闁稿�?�板畷顖炲箻椤旇棄浠掑銈嗘⒒閳峰牆顭囬妸鈺傜厓鐟滄粓宕滈悢鐓幬ュù锝囩�?�閺嬪酣鏌熼悙顒佺稇婵炲牊鍔欏娲礃閸欏鍎撳銈嗗灥濞诧箓骞嗛敓�????缁绘繈宕堕妸銏�?�闂備胶枪閺堫剟鎮疯缁綁寮�?�?顒傛崲濞戞瑦濯撮柛鎰�?级椤ユ粍銇勯妶鍜冩嫹?閿熻棄顫忕紒妯诲闁告稑锕ラ崕鎾绘⒑閻熸澘鏆辩紒缁樺浮�?�曟岸骞掗敓�????缁犲鎮归崶褍绾ф俊宸墮閳规垿鎮欓弶鎴犱户闂佹悶鍔屽﹢杈╁垝婵犳碍鏅插璺侯儑閸樹粙姊虹憴鍕凡闁告埃鍋撶紓浣靛姂椤ユ挾妲愰幒锟??惟闁靛鍠氶崥�?�攽椤旂�?�鏀绘俊鐐扮矙楠炲啴鎮滈懞銉ヤ罕闂佸壊鍋嗛崰搴ㄥ礈閸偆�???缁剧増蓱椤﹪鏌涳拷?锟筋亝鍤囬柕鍡楀暣�?�曞崬鈻庨幋鐘靛姽闁诲骸绠嶉崕閬嵥囬婊呯焼闁割偁鍨洪崰鎰扮叓閸ャ劍�???妞ゃ儲宀搁弻�???螣娓氼垱锛嗛悷婊呭鐢寮查弻銉︾厱婵炴垵宕鐐繆椤愩垼�?�伴柍瑙勫灴閸ㄩ箖宕�?懠顒勭崜婵犵绱曢崑妯煎垝濞嗗浚鍤曞┑鐘宠壘閻掓椽鏌涢幇銊︽珔妞ゅ孩鎹囧娲川婵犲啫纾╅柣蹇撶箲閻熲晛鐣烽妷褉鍋撻敐搴樺亾椤撶喐顥堥柟顔规櫊濡啫鈽夊Δ鍐╁礋闂傚�?�绀�?幗婊堝窗閹版澘绠伴柛鎰▕閸ゆ洘銇勯幇鍓佺暠缂佺姾宕电槐鎾存媴婵埈浜濈粋宥堛亹閹烘挴鎷洪梺鍛婄☉閿曪箓骞婇崘顔界厱濠电姴鍊婚崺锝忔�??閿熻姤娲樼换鍫ョ嵁鐎ｎ喗鏅搁柨鐕傛嫹?闂佽棄鍟伴崳锕傚箯閿燂拷??闂佽法鍠庨～鏇㈠磿闁�?单鍥敍濞戞﹩鍤ら梺缁橆焽缁垶鎮￠弴銏＄厸闁搞儯鍎辨俊鐓幟瑰⿰鍕闁哄本绋撻�?顒婄秵閸嬪懐浜搁幍顔剧＜缂備焦顭囩粻鎾绘煥閻曞�?�锟?????闂備胶枪椤戝懐绮旈悽鍨床婵炴垼娅曢敓锟????闂佽法鍠撻弲顐ｇ仚閻庢稒绻傞—鍐Χ閸℃浠村┑鈽嗗亝缁诲牆鐣烽崫鍕ㄦ闁靛繒濮烽娲⒑閹稿孩鈷掗柡鍜佸亰�?�曘垽宕￠悙鈺傛杸闂佺粯顭囩划顖氣槈瑜庢穱濠囶敃閿濆孩鐤佸銈冨灪濡啴骞冩禒�?�窛濠电姴瀚獮宥夋⒒娴ｅ憡鍟為柛顭戝灦閺佹捇鏁撻敓锟???????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖鎮ч崼鐔哄嚒闂佸憡鍨规慨鎾煘閹达附鍋愰悗鍦Т椤ユ繄绱撴担鍝勶拷?锟介柛銊ョ埣瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻敂閿燂拷??闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖宕滆鐢盯鏌涳拷?锟筋偓鑰块柡灞炬礋�?�曠厧鈹戦幇顓夛箓姊虹紒妯哄闁挎洩绠撻獮澶婎潰閿燂�??閿燂�??濠电偞鍨舵灙闁硅姤娲熷娲礈閹绘帊绨撮梺绋垮閻擄繝宕哄☉銏犵闁绘鏁搁敍婵囩箾鏉堝墽鍒版い顐ｇ墵椤㈡棃宕ㄩ鐓庝紟濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柡鍥ュ灩缁犲綊鎮�?☉娆樼劷闁宠棄顦甸弻宥堫檨闁告挻姘ㄩ幑銏ゅ醇閵壯冪ウ闂佸憡鍔﹂崰妤呭疾閹间焦鐓熸俊顖氭惈閺嗗崬霉濠婂嫮鐭掓慨濠冩そ�?�曟鎳栭埞鍨沪闂備礁鎼幊蹇曠矙閺嶎厼桅闁圭増婢樼粈瀣亜閺嶃劎鈻撻柟閿嬫そ濮婅櫣娑甸崨顓濇睏闂佺ǹ顑嗛惄顖氱暦濠靛鏅滃┑顔藉姃缁ㄥ姊洪棃娑辨闂傚嫬瀚悾宄扮暆鐎ｎ偄锟???闂佽法鍠曟慨銈吤哄Ο铏规殕闁归棿绀佺粻鏍喐閺傝法鏆﹀┑鍌溓归～鍛存煏韫囧﹥娅呴柡鍜佸弮濮婂宕掑▎鎴М闂佽绁撮崜婵堢箔閻旇偤鏃堝川椤撶偛浜堕梻浣虹帛閸旓箓宕滃顑芥�?�闊洦绋掗埛鎺楁煕鐏炲墽鎳呮い锔肩畵閺�?喓鍠婇崡鐐扮凹閻庡灚婢橈�??锟芥澘鐣烽崼鏇熸櫢闁跨噦�????闂佺粯甯掗悘姘跺Φ閸曨垰绠抽柛鈩冦仦婢规洜绱撴担绋库挃闁惧繐閰ｅ畷锝夊礃椤垵娈ㄩ梺瑙勫劶濡嫰鐛�?�?锛勭闁瑰鍋熼幊鍛存煕濡粯宕岄柟顔煎槻楗即宕熼鐘靛帨闁诲氦顫夊ú妯煎垝閹捐绠栭柕蹇婃濡插綊骞栧ǎ�???鐏い锟??娲栭埞鎴︽�?�鐎涙绋囬梺鍛婅壘椤戝懘鈥﹂崶褉鏋庨柟瀵稿С缁楀鈹戦悙鏉戠仧闁搞劍妞介幃锟犲即閵忋垹褰勯梺鎼炲劦椤ユ捇宕氶弶妫电懓饪伴崟顓犵厑缂備胶绮粙鎴︻敊韫囨侗鏁婇柣鎾虫捣閻嫭淇婇妶鍥ラ柛瀣洴�?�曨垶骞庨崜鍖℃�?????闂備礁鎼ú銊╁磻閹达箑纾婚柕蹇嬶�??锟介悡娆愩亜閺傛寧鎯堥柣蹇婃櫊閺岋綁鏁愯箛鏇犵槇閻庢鍠栨晶搴ㄥ箯閻樺磭鈹嶉柟鎻掝儐閿燂�???闂佽法鍠曞Λ鍕綖韫囨梻锟??婵﹩鍓涢敍婊冣攽閻愬弶顥為悽顖涘浮瀹曘垽鏁撻悩鏂ユ嫼缂備礁顑嗛娆撳磿瀹ュ鐓曢柡鍐ｅ亾闁搞劎鏁婚幃楣冩�?�閽樺宓嗛梺闈涢獜缁辨洟宕濋崼鏇燂�??锟芥鐐茬仢閸旀岸鏌熼搹顐㈠鐎殿喖顭峰畷濂稿Ψ閿�?儳骞楅梻浣虹帛閿氶柛妯荤墵閹虫粓顢旈崼鐔哄幈闂佸搫鍊搁悘婵嬵敆閵忋垻纾奸悗锝庝憾濡插憡銇勯幘鍐叉倯鐎垫澘瀚�?顒婄秵閸撴瑥顕ｉ搹顐ょ瘈闁汇垽娼ч埢鍫熺箾娴ｅ啿鍚樺☉銏╂晣闁绘劕绋勯敓锟???闁靛洦鍔欓獮鎺楀箻鐠哄搫绗氶梻鍌氾拷?锟界粈锟??鎮樺┑�?�垫晞闁告侗鍨崇粻鏃堟煙閻戞﹩娈曟い銉ユ椤潡鎳滈棃娑橆潔闂佺粯鎸堕崕鑼崲濠靛顥堟繛鎴炵懐濡倖绻濋敓�????閸曨剛顦梺璇�?�櫘閸犳牠锝炲┑瀣殝缁剧増蓱鐎氬ジ姊婚崒姘炬嫹?閿熶粙鎮ф繝鍕煓闁圭儤顧傛径濞惧牚闁割偆鍠撻崢閬嶆⒑缂佹ɑ鐓ラ柟璇х磿娴滄悂鏁傞崗鐓庮伓?闂佽法鍠撻悺鏃堝窗閺嶎叏�????閿熶粙鎮滈挊澶嬶�??锟介梺褰掑亰閸樿偐娆㈤悙娴嬫�?闁绘ɑ褰冮鎾煕閻愬瓨銇濇慨濠勭帛閹峰懘鎼归悷鎵偧闂備礁鎲″褰掞�??锟芥繝鍌ゅ殨妞ゆ劧绠戠粻鐟懊归敐鍛暈閺夊牆鐗撳娲濞戞艾顣洪梺鐟板级閿曘垹顕ｉ敓锟???瀹曞ジ鎮㈤摎鍌涚潖闂傚�?�鍊搁崐鎼佹偋婵犲嫮鐭欓柟閭�?厴閺岋附銇勮箛鎾跺闁抽攱鍨块弻鐔兼嚃閳轰椒绮舵繝纰夋嫹?閿熷鍋㈤柡�?嬬秬缁犳盯寮�?崒婊呮澖闂備浇顕栭崳锝囩不閺嶎厼绠栨繝濠傜墛鐎电姴顭跨捄铏圭伇闁哄棔鍗冲濠氬磼濞嗘垼绐楅梺鍛婄懃缁绘ê顫忔禒瀣妞ゆ牭绲鹃弲娑㈡⒑閹肩偛鍔撮柛鎾村哺閸╂盯骞掗幊銊ョ秺閺佹劙宕奸锝囩Х闂備胶枪椤戝洦绻涢埀顒勬煛鐏炲墽鈯曠紒缁樼箞瀹曟﹢顢旈崟銊ユ倕闂備胶绮幐鍫曞磹閺嶎厼绠為柕濞垮労濞撳鎮归崶顏勭处濠㈣娲栭埞鎴︽偐濞堟寧娈扮紓浣介哺濞茬喎顕ｉ銈嗗珰闁肩⒈鍓氬▓楣冩⒑缂佹ɑ鈷掗柍宄扮墦瀵偄顓奸崱妯哄伎闂佽法鍣﹂敓锟????缂佺虎鍘介幃鍌氱暦閿燂拷?鐓ゆい蹇撴噳閹风粯绻涙潏鍓ф偧闁稿簺鍊濋弫鎾绘晸閿燂拷??闂傚倷绀�?浠嬪级閸噮鐎烽梻浣烘�?缁犲秹宕硅ぐ鎺濇晣濠靛�?�枪楠炪垺绻涢崱妯曟垹绮婇鈶╂�?闁绘绮☉褔鏌涙繝鍐╋�??锟芥鐐差樀閺佹捇鎮╅崘韫暗闂備礁鎼ú銏ゅ垂濞差亝鍋傞煫鍥ㄦ惄閻斿棝鏌ら崫銉︽毄婵炴彃鐡ㄦ穱濠勭磼閵忕姵鐝濋梺璇�?�枟鏋紒鐘崇洴婵＄兘鍩￠崒銈傚亾�?�ュ鈷戦梺顐ｇ〒閳规帡鏌涢弬璺ㄐら柟骞垮灩閳规埊锟???閿熺瓔浜滅粣娑橆渻閵堝棙�???闁瑰啿绉瑰畷顐⑽旈崨顔规嫽婵炶揪绲介幉锟犲疮閻愮儤鐓熸俊銈勭贰濞堟粓鏌熼銊ユ处閸嬫劧锟???閿熻棄澹婇崰鏍�?枔閵娾晜鈷戦柛锔诲弨濡炬悂鏌ㄩ悤鍌涘�?????婵犵數濮烽弫鎼佸磻閻愬樊鐒芥繛鍡樻惄閺佸嫰鏌ㄩ悤鍌涘�???濠殿喗锚瀹曨剟寮告惔銊︾厓閻熸瑥瀚悘鎾煛娴ｅ摜效鐎规洜鍠栭�?�鏇㈠焺閸愨晝绐旈梻鍌氾�??锟介懗鑸电仚闂佹寧娲忛崕闈涚暦瑜版帒鍨傛い鏃傚亾濞堟儳鈹戦悩缁樻锭婵☆偅鐩鎶藉幢濞戞瑧鍘撻悷婊勭矒�?�曟粓鎮㈤懖鈺佺ウ闂佺鎻粻鎴︼綖閸涘瓨鐓忛柛顐ｇ箖閸ｈ姤銇勯幘铏儓妞ゎ亜鍟存俊鍫曞幢濞嗗浚娼风紓鍌欑椤戝棝宕归崸妤佹櫢闁跨噦�???????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏妞ゆ洝绮鹃ˇ褰掓煛閿燂拷?閸犳牕顫忛懡銈咁棜閻庯綆浜滅敮顖炴煟鎼淬値娼愰柟鍝ュ厴閹偤鏁傞悾灞告敵婵犵數濮村ù鍌炲极瀹ュ棛锟??闂傚牊绋掗ˉ娆愭叏鐟欏嫷娈樼紒杈ㄥ浮閹瑩顢楅�?顒勫礉閵堝鐓曟慨姗嗗墻閸庢劗绱掑畝鍐摵缂佺粯绻堝畷鍫曟嚋閸偅鐝梻鍌欒兌缁垶宕濋弴銏″仱闁靛ň鏅涘Ч鏌ユ煟濡偐甯涢柣鎾跺枛楠炴牕菐閿燂�??閻忓崬顭跨憴鍕讹�??锟介柡灞炬礋瀹曞ジ鍩楃捄铏圭Ш闁挎繄鍋犵粻娑㈠即閻樼绱叉繝纰樻閸ㄧ敻顢氳椤㈡捇骞�?崜浣猴紳婵炶揪绲芥竟濠囧磿閹扮増鍊电紒妤佺☉濞层倗澹曠憴鍕╀簻闁哄秲鍔庨妴鎺旂磼閻樿崵鐣洪柟顔筋殔閳藉鈻庡Ο鐓庡Ш闂備焦妞块崢鐓幬涘☉姘潟闁圭儤顨忛弫濠囨煟閿濆懏婀伴柛锛卞洦鈷戝ù鍏肩懅閹ジ鏌涜箛鏂嗩亪顢氶敐澶婄妞ゆ梻鈷堝濠囨⒑缂佹﹩鐒介柡浣呵归�?�鍥ㄥ緞閹邦厸鎷绘繛杈剧悼鏋い銉ョ箻閺屾冻�????閿熺瓔浜濋崳浠嬫煙楠炲灝鐏诧�??锟芥洜鍠栭�?�娑㈡晲閸℃ɑ鐝濋梻鍌欑閹诧紕鎹㈤崒婧惧亾閿燂拷?閸パ呭摋婵炲濮撮鍡涙偂閻斿憡鍙忔俊銈傚亾婵☆偅顨婂绋库槈閵忥紕鍘介棅顐㈡祫缁茶偐鑺遍悾�???纾奸弶鍫涘妼缁椦囨煙妞嬪骸鈻堟鐐存崌楠炴帡骞橀幖顓炴暢婵犵绱曢崑鎴﹀磹閵堝棛顩叉繝濠傜墕閻ゎ喗銇勯弽銊х煂闁活厼顦甸弻鐔兼倻濡崵鍘搁梺绋款儐閹瑰洭寮幇顓熷劅婵犻潧鐗婇弲濂告⒒娴ｉ涓茬紒鍙夊劤椤啴鎸婃径妯荤稁濠电偛妯婃禍婵嬎夐崼鐔虹闁瑰鍋為惃鎴︽煟閵堝懎顏慨濠呮缁瑩宕犻埄鍐╂毎闂備胶绮�?�鍫熸叏閹绢喗鍋╅柣鎴ｆ缁狅綁鏌ㄩ悤鍌涘?缂佺偓鍎抽妶鎼佸蓟閿濆绠涙い鏍ㄦ皑濮ｃ垹顪冮妶鍡樷拹闁告梹娲熼崺鐐哄箣閿旀枻锟???閿熶粙鏌涢妷銏℃珖閺嶏繝姊绘担鍛婂暈闁圭ǹ顭烽幃鐑藉煛閸涱厾鐣洪梺璺ㄥ櫐閿燂拷??濡炪們鍨哄畝鎼佸春閳ь剚銇勯幒鎴濐仼闁藉啰鍠撻�?�???绠嶉崕閬嶆偋濠婂喚鐎堕柕濞炬櫆閳锋垿鏌涘☉姗堟敾闁诡垰鐗忕槐鎺楁偐閾忣偄纰嶉梺浼欑到閸㈡煡銈导鏉戦唶闁绘棁娓圭花璇测攽閻樼粯娑ч柛濠冩�?�钘濋柟娈垮枤锟??濠囧箹缁顎嗛敓锟???娴犲鐓熼柟閭﹀墮缁狙囨煃缂佹ɑ锟??闂囧绻濇繝鍌氼�?缂佺姷鍋熼埀顒冾潐濞叉﹢宕归崸锟??鏋侀柟鍓х帛閸嬫劧�????閿熻姤娲栧ú銈夌嵁閹邦兘鏀介柣姗嗗枛閻忚鲸绻涙径�?�创闁轰礁鍟撮弫鎾绘晸閿燂�???濡炪値鍋呯换鍫熶繆閹间礁鐓涢柛灞剧矊楠炲秶绱撻崒娆戭槮妞ゆ垵鎳橀幃妯衡攽鐎ｎ亝杈堥梺缁樻濞咃絿澹曟總绋跨骇闁割偅绋戞俊浠嬫倶韫囨柨顥嬬紒杈ㄥ笒铻栭柛鎰╁妽閻忓牓鎮楃憴鍕闁稿骸銈歌棟闁规儼濮ら悡鐔哥節閸偄濮囨繛鍛У閹便劍绻濋崘鈹夸虎濡ょ姷鍋為悧鐘诲箖濞嗘挸绠甸柟鐑樼箖缂嶅�?�鈹戦悩鍨毄闁稿鐩棟濞寸厧鐡ㄩ崕搴€亜閺嶎偄鍓抽柟鍑ゆ�??闂佽法鍠曞Λ鍕綖濠靛鍤嬮柛顭戝亝閻濆啿鈹戦悩顔肩伇婵炲鐩弫鍐Ω閳轰胶顔戦梺鍝勬储閸ㄦ椽鍩涢幋锔解拻闁割偆鍠嶇欢杈ㄤ繆閹绘帞鍩ｉ柡灞剧⊕閹棃锟??閻橆偅鐏嗘俊鐐�??锟介崹娲偡閳哄懐宓�?柛銉墻閺佸洭鏌ｅΟ娲诲晱闁哥喎閰ｅ娲传閸曞灚笑闂佺粯顨呭Λ娆撳疾閸洘鍋╅敓锟???閳ь剟鎯岄幘娣簻闁瑰搫绉瑰宄懊瑰⿰鍕煁闁靛洤瀚伴獮鍥�?煛娴ｅ搫濮舵繝纰夋嫹?閿熻棄绾ч柟顔硷拷?锟藉璇差吋閸ャ劌鐝伴梺鑲┾拡閸庣柉顦查柍瑙勫灴椤㈡瑩鎮锋０浣割棜闂傚�?�鍊风欢姘焽瑜旈幃褔宕卞銏＄☉閻ｆ繈宕熼銈庡數婵犵數鍋涘Ο濠冪濠靛鍋傞柣鏂垮悑閻撶喐淇婇姘儓閻㈩垳锟??閺屻倝宕滈煫顓㈠仐闂佸搫鏈惄顖氼嚕椤掑嫭鍤勬い鏍ㄥ嚬娴煎啴姊绘担鍝ユ�?�妞ゆ泦鍛煋鐟滅増甯炲畵锟??鏌涢妷顔煎闁稿顑夐弻娑㈩敃閻樿尙浠煎Δ鐘靛仜缁夌懓顫忕紒妯诲�?�闁告稑锕ら弳鍫ユ⒑閸撹尙鍘涢柛銊ㄦ硾閻ｇ兘骞囬弶鍨敤濡炪倖鍔楅崰搴㈢閻愵剚鍙忔俊顖滃帶娴滈箖鏌ㄩ悤鍌涘�????**********************
    wire BPU_flush;
    wire inst_rreq;
    wire [31:0] inst_addr1;
    wire [31:0] inst_addr2;
    wire [31:0] BPU_pred_addr;
    wire pi_is_exception;
    wire [6:0] pi_exception_cause; 

    wire icache_inst_valid1;
    wire icache_inst_valid2;
    wire [31:0] pred_addr1_for_buffer;
    wire [31:0] pred_addr2_for_buffer;
    wire [1:0] pred_taken_for_buffer;
    wire pi_icache_is_exception1;
    wire pi_icache_is_exception2;
    wire [6:0] pi_icache_exception_cause1;
    wire [6:0] pi_icache_exception_cause2;
    wire pc_suspend;
    wire [31:0] icache_pc1;
    wire [31:0] icache_pc2;
    wire [31:0] icache_inst1;
    wire [31:0] icache_inst2;
    //*************************************************


    // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁诡垎鍐ｆ寖闂佺娅曢幑鍥灳閿燂拷?????婵＄偑鍊曠换鎰板箠韫囨挾鏆﹂柟鎯板Г閳锋垶绻涢懠棰濆殭妤犵偞鐗楁穱濠囶敃閿濆洨鐤勯悗娈垮枛椤攱淇婇幖浣哥厸闁稿本鐭花浠嬫⒒娴ｅ懙褰掑嫉椤掑倻鐭欓柟杈惧瘜閿燂拷???婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙稑鈹戦悙鏉戠亶闁瑰磭鍋ゅ畷鍫曨敆娴ｉ晲缂撶紓鍌欑椤戝棴�????閿熺獤鍥拷?锟芥い鎺戝閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁悗瑙勬礃閸ㄥ潡鐛崶顒佸亱闁割偁鍨归獮妯肩磽娴ｅ搫浜炬繝銏∶悾鐑筋敆娴ｈ鐝锋繝鐢靛У绾板秹鎮￠弴銏＄厽闁归偊鍨伴惃娲煕閳哄绋婚柟渚垮妽缁绘繈宕熼鐐殿偧闂備胶鎳撻崲鏌ュ箠濡櫣鏆﹂柕濠忓閿燂�??闂佺ǹ鏈粙鎺楁偩閼测晝纾介柛灞捐壘閳ь剟顥撶划鍫熺瑹閳ь剟鐛�?弽顓ф晝闁靛繆鏅濋崝鐑芥⒑閻愯棄鍔氱痪缁㈠弮�?�娊鏁冮崒娑氬幐闂佹悶鍎崕閬嶆�?�閳哄啰纾奸柣娆屽亾闁革綇缍佸濠氬Χ婢跺﹦鐣抽梺鍦劋閸ㄥ灚鎱ㄦ惔銊︹拺闁告稑锕ョ亸顓犵磽�?�ュ拑宸ユい顐㈢箻閹煎湱鎲撮崟顐ｏ拷?锟介梻浣告啞濞诧箓宕戦崱娴板洭濡搁埡鍌楁嫼缂備緡鍨卞ú妯衡枍閸℃稒鐓熸俊銈呭暙瀛濋梺浼欑秮�???鎲嬫�??閿熻棄銈稿鍫曞箣閻樺灚婢戦梻鍌欒兌缁垶銆冮崨瀛樺亱闊洦绋戦崒銊╂煢濡警妲撮敓�????娴犲绠抽柟鎯版绾惧綊鏌熼悧鍫熺凡缁炬儳顭烽弻鐔煎礈瑜忕敮娑㈡煟閹捐泛鏋戝ǎ鍥э躬婵�?�爼宕掑顐㈩棜濠电姷顣藉Σ鍛村磻閸涱垳鐭欓柟鎹愵嚙锟??鍡涙煙閻戞﹩娈㈤柡浣告喘閺屾洝绠涢弴鐐愩儲銇勯弬鍖�?�伐闁宠鍨堕獮濠囨煕婵犲啯宕岄柟铏殜瀹曞ジ寮撮悙鎻掍憾闂備礁缍婂Λ鍧楁倿閿曞�?�鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏缍�?弫鎾绘晸閿燂�???濠电偞鍨崹娲偂濞戙垺鐓曟繛鎴濆船閺嬨倗绱掗悩鎰佺劷缂佽鲸甯￠、姘跺幢濞嗘嚩婊堟�?�濞堝灝娅橀柛锝忕到閻ｉ攱绺介崨濠備簻闂佸憡绻傦�??锟筋剛绮绘导瀛樷拺閻犲洦鐓￠妤呮煕濡崵鐭掞拷?锟芥洘鍨块獮妯肩磼濡厧甯楅柣鐔哥矋缁挸鐣峰⿰鍫熷亜濡炲瀛╁▓鐐箾閺夋垵鎮戞繛鍏肩懇閺佹捇鏁撻敓锟????濠碉紕鍋戦崐鏍箰閻愵剚鍙忛悗闈涙憸閻牓鏌ㄩ弴鐑囨�??閿熶粙鍩涢幋鐘垫／妞ゆ挾鍋為崳铏规喐閹跺﹤鎳愮壕濂告煟濡搫鏆遍柣蹇婃櫇缁辨帡顢欏▎鎯ф闂佸疇妫勯ˇ鍨叏閳ь剟鏌ㄩ悤鍌涘?闂佺懓鍢查�?�宄邦潖濞差亜绀堥柟缁樺笂缁ㄤ粙姊洪崫銉バｉ柟鐟版喘瀹曠儤绻濋崶褍宓嗛梺缁樻⒒缁绘繄鑺辨繝姘拺闁告繂�?��?顒佹倐閹ê鈹戯拷?锟藉灚鏅滃銈嗗姂閸婃澹曟總绋跨骇闁割偅绋戞俊鏂ゆ�??閿熻姤娲栭惌澶愬箯閿燂拷??闂佽法鍠曟慨銈吤哄Ο鍏兼殰闁圭儤顨呴悡婵嬪箹濞ｎ剙濡肩紒鐘烘珪缁绘繈妫冨☉娆樻！闂佸搫妫崣鍐潖婵犳艾纾兼繛鍡樺笒閿燂拷??濠碉紕鍋戦崐鏍垂闂堟党娑樷攽鐎ｎ剙绁﹂梺纭呮彧缁犳垿鎮欓敓�??????闂備浇妫勯崯浼村窗閹邦喗宕叉繛鎴欏灩缁狅絾绻涢崱妤冪闁告梹鎸冲鐑樻姜閹殿噮妲�?梺鍝ュ枑閹稿啿顕ｆ繝姘櫜闁告稑鍊婚崰鎾诲箯閻樼粯鍤戞い鎺戯�??锟介崑鈩冪節閻㈤潧校妞ゆ梹鐗犲畷鏉课旈埀顒傚弲闂佺粯鏌ㄩ〃搴☆焽閺嶎厽鐓ｉ煫鍥ㄦ尰鐠愶紕鐥幆褍鎮戝ǎ鍥э躬椤㈡稑鈹戦幇顒侇唲闂傚�?�鍊搁ˇ顖滅矓閹绢喖鐓�?柟杈鹃檮閸婄兘鏌熺紒妯虹濡ょ姴娲ㄧ槐鎾寸瑹閸パ勭亶闂佸湱鎳撳ú顓㈠箖娴兼惌鏁婇柦妯侯槺缁愮偤姊鸿ぐ鎺戜喊闁告挻鐟х划锝呪槈濞嗘垹鐦堥梺姹囧灲濞佳冪摥闂備礁鎽滈崳銉╁磻婵犲倻鏆︽繝闈涱儏�?�告繈鎮�?☉娅辨岸骞忓ú顏呪拻闁稿本姘ㄦ晶娑氱磼鐎ｎ亞澧涢柟顖涙⒐椤︾増鎯旈敐鍥风床闂備礁鎲￠悷銉┧囨导鏉懳︽繝鍨尰閿燂拷??闂佽法鍠曟慨銈吤洪敓�????瀹曞綊宕稿Δ鍐ㄧウ濠碘槅鍨伴崥瀣舵�??閿熻姤宀搁弻銈囧枈閸楃偛鈷掑┑陇灏欐晶妤佺┍婵犲洦鍊锋い蹇撳閿燂拷??闂佽法鍠曞Λ鍕綖韫囨梻锟??婵﹩鍓欓崑宥夋偡濠婂嫭顥堟鐐诧躬楠炴鎷犻幓鎺炴�??閿熻棄顪冮妶鍡橆梿妞ゎ偄顦甸弫鎾绘晸閿燂�???闂傚倸鍊风粈�???鎮块崶顬盯宕熼�?�☉铻栭柛娑卞枛閳ь剙鐖奸弻銊モ攽閸�?晜效闂佺粯鎸搁崰娑㈠箯閿燂拷??闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍘界粩鐔煎幢濡粯鐝烽梺鍝勬储閸ㄦ椽宕戦崒鐐寸厪闁割偅绻嶅Σ褰掓煟閹惧鎳囨慨濠傤煼瀹曟帒顫濋悡搴㈩�?闂備礁鎲￠弻銊х矓瑜版帒钃燂拷?锟姐儱顦伴悡銉╂倵閿濆簼绨藉ù鐓庤嫰閳规垿顢欑涵宄颁紣濡炪値鍘奸崲鏌ユ偩闁垮闄勯柛娑橈工娴滄粓姊虹拠鈥冲箺鐎圭ǹ顭峰畷鎴﹀箻鐠囪尙顔婇梺瑙勬儗閸橀箖宕悽鍛婂仭婵犲﹤鍟撮妤呮偂閿燂�????濠电姷顣槐鏇㈠极鐠囪尙鏆﹂柣鏃傗拡閺佸秵绻涢幋鐐垫噭闁绘繃娲熷缁樻媴缁嬫妫岄梺缁樻尭閻楁挸鐣锋导鏉戝唨妞ゆ劑鍊楅敓�??????婵犳鍠栭敃銊モ枍閿濆绠柣妯款嚙閻忔娊鏌ц箛锝呬簽濞存粍鍔欏缁樼瑹婵犲啫�????闂佽法鍠曞Λ鍕嚐椤栨稒娅犳い鏍仦閻撴盯鎮楅敐搴濈暗闁稿鍨婚埀顒侇問閸犳牠骞夐敓鐘茬畾闁哄啫鐗嗘儫閻熸粌绉烽妵鎰板礋椤栨稈鎷洪梺纭呭亹閸嬫盯宕濋敂濮愪簻闁靛闄勭亸鐢电磼椤旂晫鎳勭紒缁樼箓椤繈顢橀妸锟??�????闂佽法鍠嶇划娆忣潖婵犳艾閱囬柣锟??浜介�?顒佸浮閺岋綁骞掗幘杈炬嫹?閿熶粙鏌＄仦绯曞亾�?�曞洦娈曢柣搴秵閸撴稖鎽梻鍌欐祰椤曟牠宕归崡鐐嶆盯宕�?琛″亾娴ｇ硶妲堟俊顖氬槻閻楁岸姊洪崨濠勨槈闁归攱鍨瑰濠囧礈瑜庨敓�????????婵犵妲呴崹鐢稿磻閹扮増鍋傞柣妯虹－缁犻箖鎮�?☉娆樼劷闁活厹鍊曢湁婵犲﹤绨奸柇顖氣攽閳ュ磭鎽犵紒妤嬫嫹?婵°�?�濮烽崑鐐烘晪濡炪�?�鍘煎鈥崇暦閻旂⒈鏁嗗〒姘处椤ュ牓鏌ｆ惔銈庢綈婵炴彃绻樺畷婵嬪箣閿旇�?鍋撴担绯曟�?�闁规儳纾悾楣冩偡濠婂啰肖缂侇喖顭烽幃娆徝癸拷?锟筋偅鏉搁梻浣虹帛钃辨い�???鐗犲鎶筋敍濞戞绠氶梺鍦帛鐢宕甸崶鈹惧亾鐟欏嫭绀堥柟铏崌閹�?箖鎮滈挊澶岋�??锟介悷婊冪Ч閹ɑ绻濋崒銈嗗瘜闂�?潧鐗嗗Λ娑欐櫠椤掑倻纾兼い鏃囧亹婢э箓鏌熼鎯т沪缂佺粯绻堝畷鍫曞Ω瑜嶅鎶芥⒒娴ｅ憡鎯堟繛灞傚姂�?�曟垵鈽夐姀鐘靛姦闂佽法鍣﹂敓锟????缂傚倸绉撮敃顏堢嵁閸愵喖鐏抽柡鍌樺劜椤秹鏌ㄩ悤鍌涘�??????闂傚倸鍊烽懗鍓佸垝椤栫偛�?夋俊銈傚亾闁宠绉规俊鐤槼闁哥姴妫濋弻娑㈠即閵娿儱顫梺缁樼箘閸忔ê顫忓ú顏勪紶闁告洦鍣鍫曟⒑缁嬪灝顒㈤柣鎿勭�?楠炲啴鍨鹃弬銉︼�??锟介梺鐟扮摠閺屻劍绂嶆ィ鍐╃厽闁绘柨鎲＄欢鍙夈亜韫囷絽浜滄い顓�?�劵椤﹁櫕銇勯妸銉伐闁伙絿鍏橀幖褰掝敃閵堝孩绁梺璇插嚱缂嶅棝宕戦崱娑樺偍闁汇垹鎲￠埛鎴︽煕濞戞﹫鍔熼柟鍐插暞閵囧嫰鏁傞挊澶樻婵炲瓨绮嶉幃鍌炲极閸岀偞鐓ユい鏍ㄧ煯婢规洟鏌ｉ悢鍝ユ噧閻庢凹鍘剧划鍫ュ醇閵夛妇鍘遍梺缁樏壕顓熸櫠閿燂�?????闂傚倷绀�?幖顐⒚洪�?銈呭瀭闁荤喓澧楃痪顖炴⒒閸屾埃鐪嬮柛瀣鐓ら柨鏇楀亾閻撱�?�鏌″搴�?�笧闁搞儺鍓欓悡娑㈡煕濞戝崬鏋撻柟宄邦煼濮婅櫣绮欓幐搴㈡嫳闂佽崵鍣︽俊鍥╁垝婵犲洦鍋嬮柛顐ｇ◥缁ㄥ姊洪崫鍕悙婵☆偅顨婇獮濠冨緞閹邦剛锛涢梺鍦亾閺嬬厧危閸儲鐓欓柣鎴炆戠亸浼存煟濠靛洩澹樻い顏勫暣婵�?�爼宕橀妸褌鐥梻浣藉吹閸熷潡寮插☉銏╂晪闁挎繂妫涢々鐑芥�?�閿濆懐浠涢柡鍜冪秮濮婅櫣绱掑Ο鍝勵潕闂佺ǹ绨洪崐婵嬪极瀹ュ憘鏃堝川椤旇�?�藉┑鐐舵彧閿燂�??濠殿喓鍊�?☉鐢稿醇閺囩喓鍘遍梺鎸庣箓缁绘帡鎮鹃崹顐闁绘劘灏欑粻濠氭煥閻曞�?�锟?????闂傚倸鍊峰ù鍥敋瑜嶉～婵嬫晝閸岋妇绋忔繝銏ｆ硾閳洟宕崟搴ｅ枛閹剝鎯旈敍鍕枈闂傚�?�娴囬～澶婄暦閿燂拷?椤㈡俺顦寸紒顔碱煼�?�粙顢�?悢鍝勫妇闂佽法鍣﹂敓�?????????闂傚倷鐒︽繛濠囧绩闁�?秴绀夋繛鍡樻尭閽冪喖鏌ｉ弬鍨�?�闁绘帊绮欓弫鎾绘晸閿燂�????闂備礁鎼鍐磹濠靛钃熼柨婵嗩槹閺呮彃顭跨捄铏圭伇闁哄棭鍋勯埞鎴︻敊绾嘲濮涚紓渚囧櫘閸ㄥ爼鐛箛娑樺窛妞ゆ牗绮庨悡鎾斥攽閻愬弶顥犻柛�?�崌钘熼柟杈鹃檮閳锋帒霉閿濆懏鍤堢憸鐗堝俯閺佸嫰鏌涘☉娆愮稇缂佺姷�???楠炴牗娼忛崜褍鍩岄悗娈垮枟閻擄拷?锟筋潖缂佹ɑ濯撮柛娑橈攻閸庢挾绱撴担鍓插剮缂佽埖鑹鹃悾鐑藉閵堝懐鐣鹃悷婊冪箻瀵娊濡堕崨顐熷亾閹烘埈娼╅柨婵嗘噸婢规洟姊绘担鍛婃儓闁哄牜鍓欑叅婵犻潧鐗忔稉宥嗙箾閹寸偟鎳呯紒鐘荤畺閺�?喖顢涢崱妤嬫�??閿熶粙藟濮樿埖鈷掑ù锝堟娴滃綊鏌嶅畡鎵ⅵ鐎规洘绮岄埥澶愬閳ュ厖鎮ｅ┑掳鍊х徊浠嬪疮椤栫偛鐓曢柟鐑樺灟閳ь剚甯掗～婵嬫晲閸涱剙顥氬┑鐘垫暩閸嬫﹢宕犻悩璇茬倞闁靛ǹ鍎扮純鏇㈡⒒娴ｈ櫣銆婇柛鎾寸箘缁瑩骞嬮悩鍏哥瑝濡炪�?�鐗滈崑鐐烘偂濞嗘挻鍊垫繛鎴炵懐閻掔晫绱掗悩顔煎姕缂佺粯鐩畷妤呮嚃閳轰緡娼峰┑鐑囩到濞层�?�鏁冮鍛箚闁割偅娲栧婵囥亜閹捐泛鏋戞い鏂跨Ф缁辨挻鎷呴崫鍕闂佺ǹ�?�╂繛濠冧繆閸洖绠瑰ù锝嗙摃閹芥洟姊虹紒妯烩拻闁告鍛笉闁汇垹鎲￠悡娆撴煟閹寸儐鐒界紒鐘虫崌閺屾盯骞橀弶鎴�?灆濠殿喖锕﹂崕銈忔嫹?閿熺晫鍘ч埢搴ㄥ箣濠靛棛鍘掗梻鍌欐祰椤曆呮崲閹存繄鏆嗛柟闂磋兌瀹撲線鏌涢鐘插姎閹喖姊洪幐搴㈢叆濠⒀傜矙閹線宕奸妷锔规嫼闂佸憡绋戦敃銈嗘叏閳ь剟姊洪崫鍕舵嫹?閿熶粙宕愰崷顓犵焿闁圭儤顨呴～鍛存煏閸繃顥戦柟閿嬫そ濮婃椽妫冮埡浣烘В闂佸憡鐟ラ柊锝呯暦濠靛棌鍫柛娑卞灣閿涙粎绱撻崒娆戝妽妞ゎ厼娲ㄧ划濠氬�?椤儱閰ｅ畷鎯邦檪闂婎剦鍓涢�?顒冾潐濞叉牠濡剁粙娆惧殨闁圭虎鍠楅崐鐑芥煠绾板崬澧帮�??锟芥洘妞藉濠氬磼濞嗘埈妲梺瑙勭ゴ閸撴繄绮悢鑲烘棃宕ㄩ鐙呯幢闂備礁鎲�?�ú锕傚垂闁秴纾归柤鍝ュ仯娴滄粓鐓崶銊�?鞍妞ゃ儳濮烽�?顏堝箲閹邦兛姹楃紓浣介哺閹稿骞忛崨顖涘珰闁挎稑瀚慨娲⒒閿燂�??濞佳兾涘▎鎴炴殰闁跨喓濮撮拑鐔兼煟閺傚灝顥忔俊鎻掔秺楠炴牜鍒掗悷閭﹀殥濡炪�?�甯婇梽宥嗙濠婂牊鐓ラ柡鍐ㄦ搐琚氶柣蹇撻獜缁犳捇寮婚垾宕囨殕閻庯綆鍓涜ⅵ闂備浇妗ㄩ悞锕傚礉濞嗗繒鏆﹂柕濞炬櫓閺佸秵绻涢崱妯虹伌闁崇懓绻愰埞鎴︽晬閸曨偂鏉梺绋匡攻閸ㄥ灝鐣峰┑鍥╃瘈闁搞儜鍜冪吹闂備焦鐪归崹缁樼仚缂備胶濮甸悧妤冩崲濞戙垹骞㈡俊顖濐嚙绾板秶绱撴担鍝勭彙闁搞儯鍔庨崢鐢告煟鎼淬垻鈯曟い顓炴川缁濡烽敂鍓ь啎闂佺ǹ绻楅崑鎰帮�??锟介幓鎹涘酣宕惰闊剙鈹戦垾宕囧煟鐎规洖鐖奸垾鏍敊閸濆嫬濮﹂梺鍝勬湰閸愬骞忛敓�?????闂佽法鍠撻悺鏃堝磻閸℃娲箻椤旂晫鍘搁柣蹇曞仦閺嬪鐓鍕厸濞达絿鎳撴慨鍫嫹?閿熻姤婢橈拷?锟筋厾鎹㈠┑瀣闂傚牊绋掗弳顏勨攽閻樺灚鏆╁┑顔惧厴�?�偊宕ㄦ繝鍐ㄥ伎闂佸湱铏庨崰鏍偪椤斿浜滈柟鎵虫櫅閳ь剚鐗犻�?�鏇熺鐎ｎ偆鍘介梺褰掑亰閸犳牠宕濓�??锟筋喗鐓曞┑鐘插閺嗩剟鏌＄仦璇插闁宠鍨垮畷鍗炩槈閾忣偄�????闂佽法鍠嶇划娆撳蓟濞戞鐔虹磼濡搫�?梺璺ㄥ櫐閿燂拷??????婵＄偑鍊栭崝褏寰婇悾灞筋棜闁告劕妯婂〒濠氭煏閸繂鏆欓柣蹇ｄ簼閵囧嫰濡搁妷顖氫紣闂佷紮绲块崗�???骞冮�?銏犳瀳閺夊牄鍔嶅▍鍫ユ⒒娴ｇǹ鎮戝ù�???绮欏畷鏇㈡焼瀹ュ孩鏅滈悷婊呭鐢鍩涢幒鎳ㄥ綊鏁愰崼鐕佹闂佸憡鑹剧紞濠囧蓟濞戙垺鍋愰柛鎰絻椤帡姊虹拠鈥虫灓闁稿繑锕㈤弫鎾绘晸閿燂�?????闂備胶枪椤戝棝骞愰幖渚婄稏婵犻潧顑嗛崑鍌炲箹缁顫婃繛鐓庡⒔缁辨捇宕掑▎鎴ｇ獥闂佸摜濮甸悧鐘诲箖瑜旈獮妯虹暦閸ャ劍�?????闂備胶纭堕弲婵嬪磻閻愬樊鍤楅柛鏇ㄥ灠娴肩�?鏌曟竟顖氬濞呮帡姊婚崒姘炬�??閿熶粙宕愭搴ｇ焼濞撴埃鍋撴鐐寸墵椤㈡洟鍩涘顓熴仢濠碉拷?锟界埣�?�曘劑宕掑☉姘ｆ闁剧粯鐗犻弻娑樷槈閸楃偛缁╅悶姘箖缁绘繄鍠婂Ο娲绘綉闂佽法鍣﹂敓锟??????濠电姷顣介崜婵娿亹閸愵喗鍋嬪┑鐘叉搐缁犵偤鏌曟繛鍨壔闁哄啫鐗嗛悞鐢告煥閻曞倹锟???闁捐崵鍋炵换娑㈠幢濡や胶顩伴梺鎼烇拷?锟介悧濠勬崲濞戞﹩鍟呮い鏃囧吹閸戝綊姊洪幎鑺ユ暠闁搞劌鐏濋～蹇撁洪宥嗘櫇闂�?潧鐗嗛幊宥囧垝閸洘鈷戦柛蹇撳悑閵囩喖鏌涢妸�???鎲撅�??锟筋噯锟??????缂傚倷绶￠崹鍗灻洪弽銊ь洸闁绘劦鍓涚粻楣冩煕椤愶絿绠樺ù鐘灲閺屸槄�????閿熺瓔鍋嗛埊鏇㈡煏閸パ冾伃妞ゃ垺锕㈤幃娆撳矗婢诡厸鏅涢�?�鍐Χ閸℃鈹涚紓鍌氱С缁舵岸鎮伴敓锟???閺佹捇鏁撻敓�?????濡炪們鍨洪悷褔宕版繝鍐╃秶闁靛ě鍛呯喖姊婚崒姘炬嫹?閿熶粙鎳楅崼鏇熸櫢闁跨噦�?????濠碉紕鍋戦崐鏍�?枖閿曞�?�鐐婄憸搴ㄦ倵椤掑嫭鐓熼柣鏂挎憸閹冲啴鎮�?鐓庢灓鐎殿噯锟???闂傚倸鍊烽悞锕傛儑瑜版帒鍨傞柦妯侯樈閻掔晫鎲搁弮鍫濇槬闁靛繈鍊曢柋鍥煟閺冨洦顏犳い�???娲樼换娑欐綇閸撗冨煂闂佸摜鍠庡鈥崇暦閵忋�?�绠查柟鎵虫櫃濮规姊洪崷顓炲妺闁搞劌缍婇弫宥呪堪閸愶絾�???濡炪倖娲栧Λ娑㈠礆娴煎瓨鐓曟慨姗嗗墻閸庢棃鏌熼姘伃妞ゃ垺鐩幃娆撴嚑椤掑�?�姣囧┑鐘垫暩閸嬫稑螞閿燂拷?闇夋慨妯挎硾閻ゎ噣鏌涘☉鍗炴灁濞存粍绮撻弻锟犲礃閵婏箑顦╁銈冨劚椤︾敻寮婚敐澶嬫櫆闁伙絽鐬奸悡澶娾攽椤旂�?�鍔熺紒顕呭灣缁參鎮㈤悡搴ｅ姦闂佽法鍣﹂敓�?????濡炪値鍘煎ú鈺吽囪ぐ鎺撶厵妞ゆ柣鍔屽ú銈夌嵁閵忥紕绠鹃柟瀵稿剱閻掍粙鏌ｉ妶鍛枠婵﹪缂氶妵鎰板箳閹存粌鏋堥梻浣告憸婵數鍠婂鍥╃煓濠㈣泛饪撮崥�?�煕濮樸儻�????閿熺晫绱炴繝鍥х畺闁斥晛鍟崕鐔兼煥濠靛棙顥為柛鐘崇墵濮婄粯鎷呴搹鐟扮闂佽鎮傜粻鏍х暦娴兼潙�???妞ゆ挾鍋犻幗鏇㈡⒑閻愯棄鍔氱痪缁㈠弮瀵娊濡堕崱鎰盎闂佸搫鍟ú銈夊触鐟欏嫨浜滈柨鏃囧亹閻ｉ亶妫�?敓锟?????闂備線娼荤紞鍥╃礊閿燂拷?閺佹捇鏁撻敓�???????闂備礁纾划顖炲箲閸パ呮殾鐟滅増甯╅弫濠囨煟閿濆懎顨欓梺顓у灠閳规垿鏁嶉崟顐℃�?闂佺ǹ枪閸婃繂鐣烽�?掳鍋呴柛鎰╁妿椤ρ冣攽閳藉棗鐏熼敓�????閿曞倸鍚归柡鍥╁枂娴滄粓鏌熼弶鍨暢闁伙綁浜堕弫鎾绘晸閿燂拷??闂佸憡鍔忛弬鍌涚濠婂牊鐓涢柛鎰╁妽閹兼劕霉濠婂啰绉洪柡灞剧洴�?�噣骞�?崜浣规婵＄偑鍊ゆ禍婊堝疮鐎涙ü绻嗛柛顐ｆ�?楠炪垺淇婇妶鍛殶闁瑰啿妫濆缁樻媴閸涘﹥鍠愰梺鍝ュУ閹稿寮茬捄浣曟棃宕�?鍡欏姽闁诲骸绠嶉崕閬嵥囨导瀛樻櫢闁跨噦�??????闂備緤锟???閿熻棄鑻晶鏉款熆鐟欏嫭�?冪紒鍌涘笧閳ь剨缍嗛崑鍡涘储闁�?秵鐓熼煫鍥ㄦ�?娴狅讣锟???閿熻姤娲樿摫缂佹梻鍠栭弫鎾绘晸閿燂拷??闂佸搫鑻粔鐑铰ㄩ敓�????閺屾盯骞橈拷?锟藉憡鍒涢梺璺ㄥ櫐閿燂拷????婵°�?�濮烽崑娑㈠疮閹绢喖绠栨繛鍡樻尰閸婄粯淇婇婊呭笡闁绘繃鐗犲缁樻媴閸涢潧缍婂鐢割敆閸曨�?�锔界箾閹存瑥鐏╃痪鎯ь煼閺岀喖宕滆鐢盯鏌￠崨顔剧疄闁哄本绋撴禒锕傛�?�椤掑�?�顓婚梻浣呵归敃锕傚磻濞戭澁�????閿熶粙宕�?鍢壯囨煕閳╁喚娈橀柛妯诲姉缁辨挻鎷呴崫鍕戯綁鏌涢妸褎鏆╅柛娆忔嚇濮婃椽骞愭惔銏╂闂佽桨绶￠崳锝呯暦閹达箑绠婚悗娑櫭鎾绘⒑閸涘﹤濮傞柛鏂款儏鏁堟俊銈呮噺閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曨敍濠婂懐锛滈柣搴秵閸嬪嫮绮埡鍐╁枑闁绘鐗忛惌鎺撴叏婵犲洨绱伴柕鍥ㄥ姍楠炴帡骞橈�??锟芥ɑ顔忓┑鐘殿暜缁辨洟宕戝Ο鐓庡灊婵炲棗娴氶崵鏇炩攽閻樺疇澹橀柣鎺撴そ閺屾盯骞囬埡浣割瀷缂備焦鍔楅崑銈夊蓟閿濆牏锟??闁哄洨鍋樺▽顏堟⒑閹肩偛濡界紒璇诧拷?锟介崺銏＄鐎ｅ灚鏅滈梺鍛婁緱閸ㄦ娊鎯侀崼銉︹拺闂傚牊绋撶粻鐐烘煥閻曞�?�锟?????婵犵數濮烽�?�钘壩ｉ崨鏉戠；闁告侗鍨卞畷鏌ユ煕閿燂拷?閸嬬偤宕戦埡鍐ｅ亾閻熸澘顏鐟邦儔瀵劍绂掞拷?锟筋偆鍘遍梺璺ㄥ櫐閿燂拷??闂佸搫鎳忛惄顖炵嵁閸愵喖绠ｉ柣鎰暩閻﹀牓姊洪棃娑㈢崪缂佹彃澧藉☉鐢告�?�椤戝彞绨婚梺鐟扮摠缁诲啴宕板Ο灏栧亾鐟欏嫭纾搁柛銊ょ矙楠炲啯绂掞�??锟筋亜绐涙繝鐢靛仧閸嬫搫�????閿熻棄銈稿缁樻媴閸濆嫬浠樺銈庡亝濞茬喎鐣烽幇鏉垮嵆闁靛繒濮撮崵鎴︽⒑閸濆嫸锟???閿熶粙顢栧▎鎾村亜闁糕剝鐟﹂崰鎰板箹閹碱厾鍘滈柟鍑ゆ�??闂佽法鍠曟慨銈囨崲濠靛纾兼繝濠傚椤旀洟姊绘担鍛婃儓妞わ缚鍗抽、鏍р枎韫囷絿鍔烽梺闈浥堥弲婊堟偂閺囩喆浜滈柟鎵虫櫅閳ь剚娲熷鍛婃償閳ь兛锟?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖宕滆鐢盯鏌涳拷?锟筋煉锟???閿熶粙寮婚敓鐘茬闁靛ě鍐炬毇闂傚倸鍊搁崑鍡涘垂闁�?秴桅闁告洦鍨伴崡鎶芥煥閻曞�?�锟???婵炲瓨绮撶粻鏍箖濡ゅ啯鍠嗛柛鏇ㄥ墰椤︺劑姊洪幖鐐插濠�?冮叄楠炴垿锟??閻橆偅锟??闁诲函缍嗘禍鐐哄磹閻愮儤鈷戦悗鍦У閵嗗啴鏌ら崘鑼�?煟濠碉拷?锟界埣閺佸�?�鎮鹃敓�????閻﹀牏绱掗崜褍顣奸拑杈ㄣ亜椤愵澁韬柡灞剧洴婵℃瓕顦抽柡鍡╁墰閳ь剝顫夊ú锟??宕归崸妤冨祦闁搞儺鍓﹂弫濠勭棯閹峰矂鍝烘い銉節濮婄粯鎷呴崨闈涙贡閹广垹螣娴ｆ洘绋撻幑鍕Ω閿燂拷?鎼村﹪姊虹化鏇炲⒉閼垦兠瑰⿰鍕煉闁哄矉�????閿熺瓔鍚嬮柛鎰╁妼椤�?姊哄ú璇插箹闁活厼鍊块獮鍐╃鐎ｅ灚鏅┑鐐村灦绾板秹宕氬☉銏♀拺闁告繂瀚～锕傛煕閿燂�??閸ㄥ潡鐛�?崘顔嘉у璺猴功閿涙粌鈹戦悙鏉戠仸闁挎洍鏅犻弫鎾绘晸閿燂拷????
    wire fb_pred_taken1;
    wire fb_pred_taken2;
    wire [31:0]fb_pc1;
    wire [31:0]fb_pc2;
    wire [31:0]fb_inst1;
    wire [31:0]fb_inst2;
    wire [1:0] fb_valid;
    wire [1:0]fb_pre_taken;
    
    
    wire [31:0]fb_pre_branch_addr1;
    wire [31:0]fb_pre_branch_addr2;
    wire [1:0] fb_is_exception1;
    wire [1:0] fb_is_exception2;
    wire [6:0] fb_pc_exception_cause1;
    wire [6:0] fb_pc_exception_cause2;
    wire [6:0] fb_instbuffer_exception_cause1;
    wire [6:0] fb_instbuffer_exception_cause2;

    wire [1:0]ex_is_bj;
    wire [31:0]ex_pc1;
    wire [31:0]ex_pc2;
    wire [1:0]ex_valid;
    wire [1:0]ex_real_taken;
    wire [31:0]ex_real_addr1;
    wire [31:0]ex_real_addr2;
    wire [31:0]ex_pred_addr1;
    wire [31:0]ex_pred_addr2;
    wire get_data_req;
    wire [7:0] flush_o;
    wire [7:0] pause_o;
    wire icacop_en;
    wire dcacop_en;
    wire [1:0]  cacop_mode;
    wire [31:0] cache_cacop_vaddr;

  
    wire  backend_dcache_ren;
    wire [3:0]  backend_dcache_wen;
    wire backend_dcache_writen;
    wire [31:0] backend_dcache_addr;
    wire [31:0] backend_dcache_write_data;

    // dcache 
    wire [31:0] dcache_backend_rdata;
    wire dcache_backend_rdata_valid;
    wire sc_cancel_to_backend;
    wire dcache_ready;

    // dcache-AXI 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�??????? cache 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎厽鐓㈤柛鎰典簻閺嬫盯鏌＄仦鍓ф创濠碉紕鍏橀、娆撴偂鎼搭喗娴囬梻鍌欑閹碱偊骞婅箛娑樼畺闁稿瞼鍋涢拑鐔兼煏婵炵偓娅嗛柛�?�閺佹捇鏁撻敓锟????????闂傚倸鍊搁崐鎼佸磹妞嬪海鐭嗗〒姘ｅ亾妤犵偞鐗犻�?�鏇㈡晜缂佹ɑ娅堥梻浣规偠閸庢椽宕滃▎鎴犵幓婵°倕鎳忛悡娑虫�??閿熷鍎辨鎼佺嵁閺嶎厽鐓㈤柛鎰典簻閺嬫盯鏌＄仦璇插闁诡喓鍨藉畷顐�?礋閹存瑥鐏い銊ｅ劦閹瑩顢旈崟顓濈棯濠电儑绲藉ú銈夋晝椤忓牞�????閿熻棄鈽夊Ο閿嬫杸闂佺硶鍓濆ú锟??鎯堣箛娑欌拻濞达�?娅ｇ敮娑㈡煙閸涘﹥鍊愰挊婵嬫⒒閸喍绶辨繛鍏肩墬缁绘稑顔忛鑽ょ泿婵炵鍋愰敓锟???闁哄本鐩鎾Ω閵夈儳顔掑┑鐐差嚟閸樠兠洪鐑嗘綎婵炲樊浜滄导鐘绘煏婢跺牆鍓鹃柨婵嗩槹閻撴瑩鏌涘☉姗堝伐闁告柣鍊濆畷锟犳焼�?�ュ棛鍘甸梺缁橆殔閻�?﹦娆㈤懠顒傜＜闁绘鍎ら悵顏勄庨崶褝韬┑鈥崇埣瀹曟帒顫濋銏╂婵犵绱曢崑鎴�?磹閵堝纾婚柛鏇ㄥ灠缁犵�?鏌ㄩ悤鍌涘?閻庢鍠栭�?�鐑藉极閹版澘宸濋柛灞剧矊閺嬫盯鏌熼悡搴ｇШ闁诡垰鍊垮畷顐�?Ψ瑜滃Σ绋库攽閻樺灚鏆╅柛�?�洴閹椽濡歌閸ㄦ繈鏌ｅΟ铏癸紞妞も晜鐓￠弻锝夊箛椤掑倷绮靛銈庡亝濞茬喖寮婚悢鐓庣闁�?�即娼у▓顓犵磼閻愵剙鍔ら柛姘儑閹广垹鈽夐姀鐘诧�??锟藉┑鈽嗗灥濡椼劑宕氭繝鍥ㄢ拺闁告縿鍎辨禒婊呯磽瀹ュ拑宸ユい顐㈢箻閹煎綊宕烽鐘靛幆婵犵數鍋涘Λ娆撳磿閹惰棄绀堥梺�???绉甸埛鎴︽煕閿旇骞愰柟鍑ょ�?閺屾冻锟???閿熺瓔浜烽煬顒勬煟濞戝崬鏋︾紒鐘崇☉閳藉鈻庨幇顓т户闂佽法鍣﹂敓�????????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕敐鍡╂綉闂佸搫妫旈崡鍐差潖缂佹ɑ濯撮柛娑㈡涧缂嶅﹪銆侀弽顓炲�?�婵炴垶顭囬澶愭⒑閹肩偛鍔撮柛鎾寸懇閹锋垿鎮㈤崫銉ь啎闂佺懓鐡ㄩ悷銉╂�?�閳哄懏鐓曟俊銈勭閳绘洟鏌＄仦鐐缂佺粯鐩畷褰掝敊閻撳寒娼涘┑锛勫亼閸娿�?�宕戦幒�???纾诲┑鐘插亞濞兼牗绻涘顔荤盎鐎瑰憡绻傞埞鎴︽�?�鐎靛壊鏆￠梺鎼炲妼濞硷繝鎮伴敓�????楠炲鏁冮埀顒勬倷婵犲嫭鍠愭繝濠傚枤閻掍粙鏌″搴�?�箺闁绘搫缍�?悡顐�?炊閵婏箑纰嶉柣銏╁灛閸旀垿寮诲☉姘ｅ亾閿濆骸浜濓�??锟芥洖鐬奸埀顒冾潐濞叉粓宕楅敓锟???閵嗕礁顫滈埀顒勫箖濞嗘挸绠涢柛鎾茶兌琚﹂梻浣告惈閺堫剙煤閻斿吋鏅搁柨鐕傛�????闂備礁鎼Λ�?�哥礊閿燂拷?瀵鍩勯崘鈺侊�??锟介柣鐔哥懃鐎氼剛澹曢幎鑺モ拺閺夌偞澹嗛崝宥夋煙閻熺増鍠橈拷?锟筋噮鍋婇獮妯肩磼濡粯�??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╅梻鍌ゅ灦閺屻劑寮撮悙娴嬪亾閸濄儳涓嶆い鏍仦閿燂拷????闂傚倸鍊峰ù鍥敋瑜忛�?顒佺▓閺呯娀銆佸▎鎾冲唨妞ゆ挾鍋熼悰銉╂⒑閸濆嫮鈻夐柛妯恒偢閹潡顢氶埀顒勫蓟濞戞粠妲煎銈冨妼閹虫﹢骞冮垾鏂ユ�?閻庯綆浜為鎰攽閻戝洨绉甸柛鎾寸懄娣囧﹪鎳栭埡鍐紲闂佺粯锚绾绢厼煤閹绢喗鐓涢悘鐐垫櫕鑲栭梺璇″枙閸楁娊宕规ィ鍐ㄧ闁告侗鍙庡Λ婊呯磽閸屾熬�????閿熶粙宕愰悜鑺モ挃鐎广儱顦粈澶涙嫹?閿熻В鍋撻柛鏇″煐閿燂�???闂佽法鍠曞Λ鍕偩閿熺姴绠柡鍐ｅ亾闁烩晩鍨伴悾鐑藉Ω閳轰胶顔愬銈嗘尵閸犳劕鈻嶉崶顒佲拻濞撴埃鍋撴繛浣冲懏宕查柛鈩冪☉閻掑灚銇勯幒宥囶槮濠�?屽灡娣囧﹪寮婚妷銈嗗枤濠殿喖锕︾划顖炲箯閸涱垳椹抽悗锝庡亞缁夌兘姊绘担绛嬪殐闁哥姵鐗犲畷鎰版嚒閵堝懎鐏婃繝鐢靛У閼归箖宕橀�?顒勬偡濠婂啰绠伙�??锟筋喗濞婇弫鍌炴偩閿燂拷?椤旀洟鎮楅悷鏉款棌闁哥姵娲滈懞杈ㄧ附閸涘﹦鍘搁梺鍛婁緱閸犳岸宕ｉ�?顒勬⒑閸濆嫭�?伴柣鈺婂灦�?�曟椽宕熼姘鳖槯闂佽法鍣﹂敓锟????婵炲瓨绮嶇划鎾伙�??锟藉鑸垫櫜濠㈣泛锕﹂鍥煙閼圭増褰х紒鎻掓健閹線宕奸妷锔规嫼濠殿喚鎳撳ú銈夋�?�閸欏绠惧ù锝呭暱閸熶即骞楅妷鈺傗拻闁稿本鐟ㄩ崗�?勬煙閾忣偅宕岋拷?锟芥洦鍨抽幑鍕Ω閿燂�??閿燂�????闂備線娼уΛ鏃傛濮橆剦鍤曟い鏇�?亾鐎规洖銈搁幃銏ゆ憥閸屾稓娼栫紓鍌氾�??锟介崐鎼佸磹閻戣姤鍊块柨鏇烇�??锟介�?顒婄畵�?�曞爼顢楅埀顒勫磼閵娾晜鐓熼柕蹇曞У閸熺偤鏌嶉柨�?�伌闁哄被鍊栭幈銊╁箛閼搁潧锟???闂佽法鍠嶇划娆忣嚕閹间礁绠ｉ柣鎰暩閻﹀牓姊洪棃娑氱畾婵℃彃瀚伴幊鎾诲箰鎼存稐绨婚梺闈涚箚閸撴繈藟閸喆浜滈柕蹇婃閼板潡鏌熼鐣屾噰闁糕晪绻濆畷鎺戔槈濞嗘劗甯嗛梻鍌氾�??锟介崐鐑芥�?�閿曞�?�鍑犲┑鍌溓归悿鐐箾閹存瑥鐏╅柣銈庡枟閵囧嫰寮介顫捕缂佺偓鍎崇紞濠囧蓟閻斿吋鐒介柨鏇楀亾闁告ɑ鎸抽弫鎾绘晸閿燂拷??婵炲濮撮鍡涙偂閵夛妇绠鹃柟�?�镐紳椤忓牜鏁傞柍鍝勬噺閻撴洘淇婇婊呭笡閻忓骏绠撻弻锛勪沪缁嬪灝鈷夐梺鐟板槻閹虫劗鍒掑▎鎰劅闁规儳鍘栨竟鏇㈡⒑閸撹尙鍘涢柛鐘冲哺瀵娊鏁冮崒娑氬弳濠电娀娼уΛ顓炍ｉ幖浣歌埞妞ゆ牜鍋為崑鈩冪�?婵犲倸鏆ｉ柛娆忓閳ь剚顔栭崰鏍ь嚕閸撲胶绱�?ù鐘差儏�?�告繂鈹戦悙闈涗壕閻庢矮绮欏缁樻媴閸涢潧缍婂鐢割敆閸曨剙娈炴俊銈忕到閸燁偊鎮為崹顐犱簻闁瑰搫绉堕崝宥夋煕婵犲啫濮ч柟鍑ゆ嫹?闂佽法鍠曟慨銈吤洪敓�????瀹曟繈寮介鍕喘閹囧醇閻斿嘲濡抽梻浣瑰缁诲倸煤閵娾晛绀夐悹楦匡�???�???浠嬫煟閹邦剛鎽犻悘蹇庡嵆閺屾盯鍩℃担鍛婃閻庤娲橀崹鍧楃嵁閿燂�??楠炴牠顢�?悤浣告櫖闂傚倷鑳剁划顖炲礉閺囥垺鏅搁柨鐕傛嫹???闂傚倸鍊峰ù鍥ь浖閵娾晜鍊块柨鏇烇拷?锟界粻鏌ユ煕閵夘喖澧紒鐘崇墵閺屽秹宕崟锟??娅ら梺鎼烇拷?锟介崹鍫曞Φ閸曨垰绠抽柟鎼幗绗戦梻浣芥�?�锟??浣虹礊婵犲偆娼栧┑鐘宠壘绾惧吋绻涢崱妯虹劸婵″樊鍠氱槐鎾诲磼濮樻瘷銏ゆ煥閺囨﹫锟???閿熶粙鎮橈拷?锟筋喗鐓熼柣妯哄帠閼割亪鏌涢弬鍧�?弰闁诡垰鐭傚畷鍗烆渻閺囩偟绉洪柡浣瑰姍�?�曘劑顢欓崗鍏肩暭缂傚�?�鍊烽懗鍫曟惞鎼淬劌鍨傞悹杞拌濞兼牕鈹戦悩瀹犲缁炬儳鍚嬬换娑㈠幢濡櫣鍔稿┑鈥虫▕閸犳氨妲愰幘璇茬＜婵ɑ鐦烽�?銈嗙叆闁哄洦锚閳ь剚鐩幃姗堟�??閿熺瓔鍠楅悡鐔兼煟濡搫甯犻柤鍓蹭邯閺屾盯寮崸�???寮伴梺璇″灠閻倸鐣烽崡鐑嗘富闁哄洨鍋熺粔娲煛娴ｇ懓濮嶏拷?锟芥洖銈搁幃銈嗘媴�?�勭増鎲㈠┑鐘垫暩閸嬬偤宕归崼鏇炵闁告縿鍎抽惌鎾舵喐閻�?牆绗掗柦鍐枛閺屽秹濡烽敓锟???婢ь垶鏌涘顒夊剶闁哄本鐩獮鍥煛娴ｅ壊鐎抽梺璇″灣閸犲酣鍩為幋锔斤�??锟介柤纰卞墯閹茶偐绱撴笟鍥ф灈缂佸鐖煎畷姘跺箳閿燂拷?缁犲鎮归崶顏勮敿闁硅姤娲熷铏规崉閵娿儲鐏佹繝娈垮枟閹告娊骞冨▎鎰瘈闁搞儯鍔庨崢鎾绘煛婢跺苯浠у褎顨婅棟闂佸灝顑囩粻鎾呮�??閿熻В鍋撳┑鐘辫兌閻╁骸顪冮妶搴濈盎闁哥喎鐡ㄦ穱濠囧醇閺囩偟顦ㄩ梺闈浨归崕杈暯闂傚�?�鍊烽懗鑸电仚濡炪�?�鍨甸崯鏉戠暦閹邦兘�?介悗锝庡墮缁侊箓姊洪崨濠傚闁告搩鍣ｅ�???宕煎┑鍫濆Е婵＄偑鍊栫敮鎺炴嫹?閿熻棄鎽滅槐鐐哄�?閵娧呯槇闂傚倸鐗婃笟妤呭磿閹扮増鐓曞┑鐘叉处閺侀亶鏌曢崶褍顏鐐村浮�?�曞崬顪冮幆褜妫滄繝纰夌磿閸嬫垿宕愰弴銏℃櫢闁跨噦锟??????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛锟??????闂傚倸鍊搁崐椋庣矆閿燂拷?楠炲鏁撻悩鍐蹭画闂�?潧锛忛崟顐㈢哎闂佽法鍣﹂敓锟?????闁诲孩顔栭崰鏍�??锟藉畡閭�?殨闁圭虎鍠栭～鍛存煟濡鍤欓柡浣筋潐缁绘繈鎮介棃娴躲垽鏌ｈ箛鏂垮摵鐎规洘绻堝浠嬪Ω閿旂晫褰欓梻鍌氾�??锟介崐鎼佸磹妞嬪海鐭嗗�?�姘ｅ亾妤犵偞鐗犻�?�鏇㈡晝閳ь剛绮婚鐐达拷?锟介柨婵嗛�?�娴滅偞銇勯埡浣哥骇闁靛洤�?�粻娑㈠箻閹颁椒绱濇繝鐢靛仜閸氬鎮у⿰鍛潟闁规儳鐡ㄦ刊鎾煠濞村澧查柛銊ョ埣�?�曟碍绻濋崶褏顔掑銈嗘⒒閺咁偊宕㈡ィ鍐┾拺閻犲浄锟???閿熻棄绠洪柣銏╁灡鐢拷?锟界暦濠靛围濠㈣泛顑囬崢顏堟⒑缁洖澧叉い銊﹀姍閻擃剟顢楁担鐟板伎婵犵數濮撮崯顖炲Φ濠靛洣绻嗘い鎰╁灩閺嗭綁鏌涢埡�?�瘈鐎规洘锕㈤、鎾活敍濡�?鍋撳Δ鍐╊潟闁规儳鐡ㄦ刊鎾煕濠靛棗鐝旈柨婵嗩槹閻撴瑩鏌ｉ悢鍝勵暭闁哥姵锕㈤弻鐔碱敊鐠囨彃绁銈冨灪閻熝囧箲閸曨垰惟鐟滃骸顭块幋鐐电瘈闁汇垽娼ф禒锕傛煕閵娿儳鍩ｉ柟顔惧厴閺佹捇鏁撻敓�?????闂佸疇顕х粔瑙勬叏閳ь剟鏌曢崼婵囶棏闁归攱妞介弻锝夋偐閸忓懓鍩呴梺鍛婃煥閼活垶鍩㈠澶婄�?闁绘鐗忛崢鐢告⒑閸涘﹤鐏熼柛濠冪墵閺佹捇鏁撻敓�???????
    wire dev_rrdy_to_cache;
    wire dev_wrdy_to_cache;

    wire duncache_rvalid;
    wire [31:0] duncache_rdata;
    wire  duncache_ren;
    wire [31:0] duncache_raddr;

    wire duncache_write_finish;
    wire duncache_wen;
    wire [31:0] duncache_wdata;
    wire [31:0] duncache_waddr;
    
    wire [31:0] new_pc_from_ctrl;
    wire [1:0] BPU_pred_taken;

    //闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧懓顪冿拷?锟筋亝鎹ｉ柣顓ㄦ�???婵°�?�濮烽崑娑⑺囬悽绋挎瀬闁瑰墽绮崑鎰版煕閹邦剙绾ч柣銈呭濮婄粯鎷呯粵瀣異闂佹悶鍔岄妶鎼佸箖閿燂�??楠炲洭顢涘Ο瑙勭潖闂佽法鍣﹂敓�?????????缂傚倸鍊搁崐鐑芥倿閿斿墽鐭欓柟杈惧瘜閺佸嫰鏌涢埄鍐槈闁汇�?�鍋撶换婵囩�?閸屾碍鐏撳┑鐐存尭椤兘寮婚弴銏犻唶婵犻潧娴傚Λ鐐电磽娴ｈ娈曢悽顖ょ�?楠炲啫螖閳ь剟锝炲┑�?�亗閹艰揪绱曢惈鍕煟鎼淬値娼愭繛鍙壝叅闁哄稁鍙庨弫鍥煕韫囨洖甯剁紒鍓佸仱閹鏁愭惔鈥愁潻濡ょ姷鍋涢悧鎾愁潖缂佹ɑ濯撮柛娑橈龚閿燂�??闂備胶枪缁ㄦ椽宕愬Δ鍛闁靛繈鍊曠粈鍐煏婵炲灝鐏柣蹇ユ嫹???婵犵數鍋涘Ο濠冪濠靛鐓曢柟鐑樺殮瑜版帗鏅查柛娑卞枛閺嗗牓姊虹拠鈥崇仩闁绘锕俊鐢稿礋椤栨稒娅嗛柣鐘叉穿鐏忔瑦绂掗幖浣光拺閻犲浄锟???閿熻姤娈梺鍛婃处閸�?箖鎯�?崼銉︹拺闁硅偐鍋涢敓�????闂佸憡绮堢粈�???寮ぐ鎺撯拻闁稿本鐟чˇ锔剧磽�?�ュ拑宸ラ敓�?????????闂備浇顕栭崹浼存嚐椤栨繄浜欓梻浣告啞娓氭宕板璺哄偍闂侇剙绉甸埛鎴︽煛閸屾ê鍔滄繛鍛嚇閺屾盯鎮㈢捄鍝勭ギ濡ょ姷鍋涢敃顏勭暦閵娾晩鏁嶆繝濠傚缁憋繝姊绘担绛嬪殐闁搞劌閰ｅ畷�???鍩★�??锟筋偄锟???闂佽法鍠曟慨銈囨崲濞戙垺鏅查柛娑卞枟閹瑩姊洪幐搴㈠濞存粠浜悰锟??宕橀妸銏★拷?锟介梺鐟扮仢閸燁垶寮查姀銈嗏拺缂佸鍎婚～锕傛煕婵犲啰澧碉拷?锟筋喛灏欏濠傤潡椤хaddr闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌ｉ幋锝呅撻柛濠傛健閺屻劑寮撮悙娴嬪亾瑜版帒纾块柟瀵稿У閸犳劙鏌ｉ敓�????閻楀棛绮幒妤佹櫢闁跨噦�????????闂備緤锟???閿熻棄鑻晶鎾煥閻曞�?�锟???闂佽法鍣﹂敓�????????濠碉紕鍋戦崐鏍暜婵犲嫮鐭嗗〒姘ｅ亾鐎规洜鏁婚弫鎾绘晸閿燂拷??闂傚洤顦扮换婵囩�?閸屾凹锟??缂備胶濮甸�?�鍥╂閹烘鏁婇柣锝呯焾閺嗭拷?锟解攽閻愰潧甯剁紒缁樕戞穱濠傤潰�???濠冃梻浣风串缁犳垿鎮ч幘鎰佹綎婵炲樊浜滅粻褰掓煟閹邦厼绲诲┑鈯欏洦鈷戦柛娑橈梗缁堕亶鏌ㄩ悤鍌涘???闂傚倸鍊搁崐鎼佸磹閹间礁纾癸�??锟藉嫭鍣磋ぐ鎺戠倞鐟滃寮搁弽顓熺厸闁搞儯鍎遍悘鈺呮⒒閸屻�?�鐏﹂柡灞诲姂�?�挳鎮滈崶銊ヮ�??闂佽法鍠撻弲顐ゅ垝婵犳凹鏁嶉柣鎰嚟閸欏棝姊虹紒妯荤闁稿﹤缍婇弫鎾绘晸閿燂�???
    wire [31:0] csr_dmw0;//dmw0闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌ｉ幋锝呅撻柛濠傛健閺屻劑寮崼鐔告闂佺ǹ顑嗛幐鍓у垝椤撶偐妲堟俊顖濐嚙濞呇囨⒑濞茶骞楅柣鐔叉櫊�?�鎮㈤崨濠勭Ф闂佸憡鎸嗛崨顔筋啅闂備浇顕э拷?锟解晠鎳濇ィ鍏洦�?�奸弶鎳筹箓鏌涢弴銊ョ仩缂佺姵濞婇弻娑㈠焺閸愶缚娌繝銏ｎ潐濞茬喎顫忕紒妯诲闁荤喖鍋婇崵�?�攽閻愭潙绲荤紒缁樏悾椋庢喆閸曨収娴勯柣搴秵娴滄繈鎮楅鍕拺闁荤喐婢�?埛鏃傜磼椤曞懎鐏︼拷?锟筋喗鐓￠獮鏍ㄦ媴閸︻厼寮抽梻浣虹帛濞叉牠宕愯ぐ鎺撴櫢闁跨噦�?????闂傚倸鍊峰ù鍥敋瑜忛�?顒佺▓閺呯娀銆佸▎鎾冲唨妞ゆ挾鍋ら敓�??????闁诲氦顫夊ú锟??宕归崜浣瑰床婵犻潧顑呯壕鍏肩�?婵犲倸顏い�???娲熷缁樻媴閾忕懓绗￠梺鍦归幗婊堟嚍闁�?秴閱囬柡鍥╁仱閸炶泛顪冮妶鍛闁绘锕幃锟犲即閻旇櫣顔曢梺鐟扮摠缁诲倿鎳滆ぐ鎺撶厽閹兼番鍨洪妵婵嬫煛鐏炵偓绀夌紒鐙呮�?????闂傚倷鐒︽繛濠囧绩闁�?秴鍨傞柛褎顨呴拑鐔哥箾閹寸�?�姘跺绩娴犲鐓曢柍鈺佸枤濞堛垹霉閻�?潧甯舵い顏勫暣婵″爼宕ㄩ缁㈡炊闂備胶枪椤戝懘鏁冮鍕靛殨濠电姵鑹炬儫闂佸啿鎼崐鍛婄閻愮儤鈷戠紒瀣锟??鎵磼鐎ｎ偄鐏存い顫嫹??27:25]闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌ｉ幋锝呅撻柛濠傛健閺屻劑寮崼鐔告闂佺ǹ顑嗛幐鍓у垝椤撶偐妲堟俊顖濐嚙濞呇囨⒑濞茶骞楅柣鐔叉櫊�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戦柟鑲╁仜閳ь剚鐗犲畷婵嬪�?椤撶倣锕傛煕閺囥劌鐏犻柛鎰ㄥ亾闂備線娼ц噹闁告侗鍨抽悰銉︾�?閻㈤潧浠滈柣掳鍔庨崚鎺戠暆閳ь剛妲愰悙瀵哥瘈闁搞儜鍡樻啺闂備焦瀵х粙鎴�??閿熺瓔浜滈埢浠嬵敂閸喎浠梺鎼炲劘閸斿瞼寰婄拠娴嬫�?妞ゆ棁濮ょ粈瀣叏婵犲啯銇濇鐑囨嫹???????濠电偞娼欓崥瀣焽濞嗘挻瀚呴柣鏂垮悑閻撶喖鏌￠崘銊︾カ闁瑰嚖�?????闂備胶枪椤戝棝骞愰幖浣哥�?濠㈣泛艌閺嬪秵銇勯幘�???鍊婚弫鏍磽娓氬洤娅�?柛娆屽亾濡炪倧绠戦顓犳閹烘挻缍囬柕濞垮劜鐠囩偛螖閻橀潧浠滄繛宸弮閵嗕礁螣濞嗙偓歇闂備椒绱徊浠嬫偉閻撳寒娼栧┑鐘宠壘閻愬﹦鎲稿⿰鍫熸櫢闁跨噦锟???闂傚倷绀�?幖顐ゆ偖椤愶箑绀夐敓�????閸曨偆鍘撮梺纭呮彧缁犳垿鐛�?鈩冨弿婵°倐鍋撴俊顐ｇ懇閺佹捇濡烽埡鍌楁嫽婵炶揪锟??椤濡甸悢鍏肩厱婵☆垳鍘х敮鍫曟懚閻愬�???闂傚牊渚楅崕蹇曠磼閻樺磭澧遍柟鍙夋�?�閹囧醇濠靛牏鎳嗙紓鍌欒兌婵數绮欓幒�???桅闁告洦鍨板Λ�???鏌涢…鎴濇灍闁稿⿴鍨跺铏规嫚閼碱剛顔囬梺缁橆殕閹瑰洭鐛�?崘顔芥櫢闁跨噦锟???闂佸磭绮幑鍥х暦瑜版帩鏁婇柣锝呭婢规洟姊婚崒娆愮グ婵℃ぜ鍔庣划鍫熺瑹閳ь剟鍨鹃敓�????閻ｏ繝骞嶉鑺ヮ啎闂佽法鍣﹂敓锟???????濠碉紕鍋戦崐鏍暜婵犲洦鈷旓�??锟姐儱妫涢�?�鍙夌節婵犲倻澧涢柣鎾寸懇閺岋綁骞嬮悘娲讳邯閹﹢濡烽敂杞扮盎闂婎偄娲ら敃銉モ枍婵犲洦鐓欐い鏃傚帶濡插鏌嶇拠鏌ワ拷?锟介柍璇查叄楠炲鎮╅搹顐晫婵犲痉甯�??閿熻姤鎱ㄩ悜钘夌；闁绘劗鍎ら崑�?�煛閸ワ絺鍋撳畷鍥锋嫹?閿熻棄鈹戦敍鍕杭闁稿﹥鐗曢蹇旂節濮橆剛锛涢梺鐟板⒔缁垶鎮￠崘顏呭枑婵犲﹤鐗嗙粈鍫熸叏濡灝鐓愰柛�?�儐缁绘繃绻濋崒娑樻闂佹悶鍔嶇换鍌炲煘閹达附鍋愰柛娆忣槺閵堚晠姊烘潪鎵槮妞ゆ垵顦靛璇差吋閸偅顎囬梻浣告啞閹搁箖宕版惔顭戞晪闁挎繂妫涢敓�????濠殿喗锕╅崢鍏肩濠婂牊鈷戦柛蹇氬亹閵堟挳鏌￠崨顔撅�??锟界紒顔硷躬閺佸啴宕掑☉鎺撳闂備礁鎲￠幑浣轰焊濞嗘挸鍌ㄦ繛鎴欏灪閻撴洟鏌ｅΟ铏癸紞妞わ綀灏欑槐鎺�?磼濞戞鐟茬紓浣芥�?�缁瑥鐣烽妸锔剧闁绘劦鍓欓褰掓⒒閸屾瑨鍏屾い銏狅躬瀹曟垿骞囬弶璺紱濠电偞鍨崹褰掓�?�閻㈠憡鏅搁柨鐕傛嫹?????闂佽姘﹂～澶娒洪埡鍐濞达絽鎽滈弳锕傛煥閻曞倹锟???闂佺偨鍎荤粻鎾荤嵁鐎ｎ亖�?介柛銉ㄦ硾閹亪姊婚崒姘炬嫹?閿熺晫绮堟担鍦彾濠电姴娲ょ壕濠氭煕濞戝崬濮告繛宸簻閿燂拷?閻熸粌閰ｅ鍐测堪閸啿鎷洪梺鐓庮潟閸婃洟寮搁幋鐘电＜妞ゆ棁鍋愰悞鎼佹煛鐏炴枻韬柡浣瑰姈�?�板嫭绻濋崟顓熸瘒婵犲痉甯�??閿熺晫寰婃禒瀣柈妞ゆ牜鍋為崐鍧楁煥閻曞倹锟????濡ょ姷鍋涢悘婵嬪礉濮橆厺绻嗘い鎰剁悼濞茶揪锟???閿熻姤娲忛崹浠嬪蓟閸℃鍚嬮柛鈥崇箲鐎氬ジ姊绘担鍛婅�?閺嬵亪鎮�?☉鎺撴珚閽樼喖鏌涢埄鍐︿粶閿燂拷?娴犲鏅搁柨鐕傛�??????濠电姷鏁搁崑娑樜涙惔銊ュ瀭闁芥ê顦遍弳锕傛煥濠靛棙顥滅紒鍓佸仱閺佹捇鏁撻敓�??????婵＄偑鍊栧鐟懊洪悢濂夋綎闁惧繐�?辩壕鍏间繆椤栨繍鍤欑痪鏉跨У娣囧﹪濡堕崶顬綁鏌熼纭锋嫹?閿熶粙顢氶敐澶婄闁兼亽鍎插▍婊勭節閵忥絾纭炬い鎴濇喘�?�曘垽妫冨☉杈ㄥ瘜闂�?潧鐗嗗Λ娑欐櫠椤掑嫭鐓犵憸鐗堝笧閻ｇ尨�????閿熺瓔鍠楁繛濠囧极閹版澘鐐婇柨婵嗘噸婢规洟鏌ｉ悢鍝ユ噧閻庢凹鍘剧划鍫ュ醇閵夛妇鍘遍梺缁樏壕顓熸櫠閻㈠憡鐓忛柛鈩冩礈椤︼箓鎽堕弽顬�?�綊鏁愰崶銊ユ畬濡炪倕�?�╅幐缁樼┍婵犲洦鍊凤拷?锟藉壊鍠栭崜鐗堜繆閵堝洤孝闁硅姤绮庨崚鎺楊敇閵忕姷鍔撮梺鍛婂姦娴滅偤鎯侀崼銉︼拷?锟介柛蹇暻瑰畵鍡涙煛閳ь剟宕￠悜鍡欏數闂佽法鍣﹂敓�?????闂佽法鍣﹂敓�?????婵＄偑鍊栫敮濠囨倿閿斿墽鐭嗛悗锝堝煐閿燂�???闂佽法鍠曟慨銈吤洪敓�????瀹曟繂鈻庤箛鏇熸闂佺粯鍨归悺鏃堝极閸ヮ剚鐓熼柡鍐ㄦ处椤忕娀鏌￠崱鎰伄缂佽鲸鎹囧畷鎺戭潩閻愵剙�????闂佽法鍠嶇划娆忕暦閹扮増鍊婚柤鎭掑劚閳ь剙娼￠弻銊╁即閻愭祴鍋撻崨濠庢敯闂傚�?�鑳剁划顖炲礉濡ゅ懎纾块柕鍫濐槸绾惧綊鏌涜椤ㄥ棝鎮￠妷鈺傛櫢闁跨噦�????????缂傚倸鍊烽懗鑸靛垔椤撱垹鍨傞柛顐ｆ礀閽冪喐绻涢幋鐐冩艾危閸喍绻嗘い鏍ㄨ壘閹垿鏌熼幓鎺嬪仮婵﹥妞藉畷顐﹀礋閿燂拷?濞呫倝姊虹拠鈥虫灈闁稿﹤鐏濋锝嗙節濮橆儵鈺呮煃閸濆嫸锟???閿熻姤绂嶉悙鐑樷拺缂佸瀵у﹢鎵磼鐎ｎ偄鐏存い顫嫹??
    wire [31:0] csr_dmw1;//dmw1闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌ｉ幋锝呅撻柛濠傛健閺屻劑寮崼鐔告闂佺ǹ顑嗛幐鍓у垝椤撶偐妲堟俊顖濐嚙濞呇囨⒑濞茶骞楅柣鐔叉櫊�?�鎮㈤崨濠勭Ф闂佸憡鎸嗛崨顔筋啅闂備浇顕э拷?锟解晠鎳濇ィ鍏洦�?�奸弶鎳筹箓鏌涢弴銊ョ仩缂佺姵濞婇弻娑㈠焺閸愶缚娌繝銏ｎ潐濞茬喎顫忕紒妯诲闁荤喖鍋婇崵�?�攽閻愭潙绲荤紒缁樏悾椋庢喆閸曨収娴勯柣搴秵娴滄繈鎮楅鍕拺闁荤喐婢�?埛鏃傜磼椤曞懎鐏︼拷?锟筋喗鐓￠獮鏍ㄦ媴閸︻厼寮抽梻浣虹帛濞叉牠宕愯ぐ鎺撴櫢闁跨噦�?????闂傚倸鍊峰ù鍥敋瑜忛�?顒佺▓閺呯娀銆佸▎鎾冲唨妞ゆ挾鍋ら敓�??????闁诲氦顫夊ú锟??宕归崜浣瑰床婵犻潧顑呯壕鍏肩�?婵犲倸顏い�???娲熷缁樻媴閾忕懓绗￠梺鍦归幗婊堟嚍闁�?秴閱囬柡鍥╁仱閸炶泛顪冮妶鍛闁绘锕幃锟犲即閻旇櫣顔曢梺鐟扮摠缁诲倿鎳滆ぐ鎺撶厽閹兼番鍨洪妵婵嬫煛鐏炵偓绀夌紒鐙呮�?????闂傚倷鐒︽繛濠囧绩闁�?秴鍨傞柛褎顨呴拑鐔哥箾閹寸�?�姘跺绩娴犲鐓曢柍鈺佸枤濞堛垹霉閻�?潧甯舵い顏勫暣婵″爼宕ㄩ缁㈡炊闂備胶枪椤戝懘鏁冮鍕靛殨濠电姵鑹炬儫闂佸啿鎼崐鍛婄閻愮儤鈷戠紒瀣锟??鎵磼鐎ｎ偄鐏存い顫嫹??27:25]闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌ｉ幋锝呅撻柛濠傛健閺屻劑寮崼鐔告闂佺ǹ顑嗛幐鍓у垝椤撶偐妲堟俊顖濐嚙濞呇囨⒑濞茶骞楅柣鐔叉櫊�?�鎮㈤崨濠勭Ф婵°�?�绲介崯顖烆敁�?�ュ鈷戦柟鑲╁仜閳ь剚鐗犲畷婵嬪�?椤撶倣锕傛煕閺囥劌鐏犻柛鎰ㄥ亾闂備線娼ц噹闁告侗鍨抽悰銉︾�?閻㈤潧浠滈柣掳鍔庨崚鎺戠暆閳ь剛妲愰悙瀵哥瘈闁搞儜鍡樻啺闂備焦瀵х粙鎴�??閿熺瓔浜滈埢浠嬵敂閸喎浠梺鎼炲劘閸斿瞼寰婄拠娴嬫�?妞ゆ棁濮ょ粈瀣叏婵犲啯銇濇鐑囨嫹???????濠电偞娼欓崥瀣焽濞嗘挻瀚呴柣鏂垮悑閻撶喖鏌￠崘銊︾カ闁瑰嚖�?????闂備胶枪椤戝棝骞愰幖浣哥�?濠㈣泛艌閺嬪秵銇勯幘�???鍊婚弫鏍磽娓氬洤娅�?柛娆屽亾濡炪倧绠戦顓犳閹烘挻缍囬柕濞垮劜鐠囩偛螖閻橀潧浠滄繛宸弮閵嗕礁螣濞嗙偓歇闂備椒绱徊浠嬫偉閻撳寒娼栧┑鐘宠壘閻愬﹦鎲稿⿰鍫熸櫢闁跨噦锟???闂傚倷绀�?幖顐ゆ偖椤愶箑绀夐敓�????閸曨偆鍘撮梺纭呮彧缁犳垿鐛�?鈩冨弿婵°倐鍋撴俊顐ｇ懇閺佹捇濡烽埡鍌楁嫽婵炶揪锟??椤濡甸悢鍏肩厱婵☆垳鍘х敮鍫曟懚閻愬�???闂傚牊渚楅崕蹇曠磼閻樺磭澧遍柟鍙夋�?�閹囧醇濠靛牏鎳嗙紓鍌欒兌婵數绮欓幒�???桅闁告洦鍨板Λ�???鏌涢…鎴濇灍闁稿⿴鍨跺铏规嫚閼碱剛顔囬梺缁橆殕閹瑰洭鐛�?崘顔芥櫢闁跨噦锟???闂佸磭绮幑鍥х暦瑜版帩鏁婇柣锝呭婢规洟姊婚崒娆愮グ婵℃ぜ鍔庣划鍫熺瑹閳ь剟鍨鹃敓�????閻ｏ繝骞嶉鑺ヮ啎闂佽法鍣﹂敓锟???????濠碉紕鍋戦崐鏍暜婵犲洦鈷旓�??锟姐儱妫涢�?�鍙夌節婵犲倻澧涢柣鎾寸懇閺岋綁骞嬮悘娲讳邯閹﹢濡烽敂杞扮盎闂婎偄娲ら敃銉モ枍婵犲洦鐓欐い鏃傚帶濡插鏌嶇拠鏌ワ拷?锟介柍璇查叄楠炲鎮╅搹顐晫婵犲痉甯�??閿熻姤鎱ㄩ悜钘夌；闁绘劗鍎ら崑�?�煛閸ワ絺鍋撳畷鍥锋嫹?閿熻棄鈹戦敍鍕杭闁稿﹥鐗曢蹇旂節濮橆剛锛涢梺鐟板⒔缁垶鎮￠崘顏呭枑婵犲﹤鐗嗙粈鍫熸叏濡灝鐓愰柛�?�儐缁绘繃绻濋崒娑樻闂佹悶鍔嶇换鍌炲煘閹达附鍋愰柛娆忣槺閵堚晠姊烘潪鎵槮妞ゆ垵顦靛璇差吋閸偅顎囬梻浣告啞閹搁箖宕版惔顭戞晪闁挎繂妫涢敓�????濠殿喗锕╅崢鍏肩濠婂牊鈷戦柛蹇氬亹閵堟挳鏌￠崨顔撅�??锟界紒顔硷躬閺佸啴宕掑☉鎺撳闂備礁鎲￠幑浣轰焊濞嗘挸鍌ㄦ繛鎴欏灪閻撴洟鏌ｅΟ铏癸紞妞わ綀灏欑槐鎺�?磼濞戞鐟茬紓浣芥�?�缁瑥鐣烽妸锔剧闁绘劦鍓欓褰掓⒒閸屾瑨鍏屾い銏狅躬瀹曟垿骞囬弶璺紱濠电偞鍨崹褰掓�?�閻㈠憡鏅搁柨鐕傛嫹?????闂佽姘﹂～澶娒洪埡鍐濞达絽鎽滈弳锕傛煥閻曞倹锟???闂佺偨鍎荤粻鎾荤嵁鐎ｎ亖�?介柛銉ㄦ硾閹亪姊婚崒姘炬嫹?閿熺晫绮堟担鍦彾濠电姴娲ょ壕濠氭煕濞戝崬濮告繛宸簻閿燂拷?閻熸粌閰ｅ鍐测堪閸啿鎷洪梺鐓庮潟閸婃洟寮搁幋鐘电＜妞ゆ棁鍋愰悞鎼佹煛鐏炴枻韬柡浣瑰姈�?�板嫭绻濋崟顓熸瘒婵犲痉甯�??閿熺晫寰婃禒瀣柈妞ゆ牜鍋為崐鍧楁煥閻曞倹锟????濡ょ姷鍋涢悘婵嬪礉濮橆厺绻嗘い鎰剁悼濞茶揪锟???閿熻姤娲忛崹浠嬪蓟閸℃鍚嬮柛鈥崇箲鐎氬ジ姊绘担鍛婅�?閺嬵亪鎮�?☉鎺撴珚閽樼喖鏌涢埄鍐︿粶閿燂拷?娴犲鏅搁柨鐕傛�??????濠电姷鏁搁崑娑樜涙惔銊ュ瀭闁芥ê顦遍弳锕傛煥濠靛棙顥滅紒鍓佸仱閺佹捇鏁撻敓�??????婵＄偑鍊栧鐟懊洪悢濂夋綎闁惧繐�?辩壕鍏间繆椤栨繍鍤欑痪鏉跨У娣囧﹪濡堕崶顬綁鏌熼纭锋嫹?閿熶粙顢氶敐澶婄闁兼亽鍎插▍婊勭節閵忥絾纭炬い鎴濇喘�?�曘垽妫冨☉杈ㄥ瘜闂�?潧鐗嗗Λ娑欐櫠椤掑嫭鐓犵憸鐗堝笧閻ｇ尨�????閿熺瓔鍠楁繛濠囧极閹版澘鐐婇柨婵嗘噸婢规洟鏌ｉ悢鍝ユ噧閻庢凹鍘剧划鍫ュ醇閵夛妇鍘遍梺缁樏壕顓熸櫠閻㈠憡鐓忛柛鈩冩礈椤︼箓鎽堕弽顬�?�綊鏁愰崶銊ユ畬濡炪倕�?�╅幐缁樼┍婵犲洦鍊凤拷?锟藉壊鍠栭崜鐗堜繆閵堝洤孝闁硅姤绮庨崚鎺楊敇閵忕姷鍔撮梺鍛婂姦娴滅偤鎯侀崼銉︼拷?锟介柛蹇暻瑰畵鍡涙煛閳ь剟宕￠悜鍡欏數闂佽法鍣﹂敓�?????闂佽法鍣﹂敓�?????婵＄偑鍊栫敮濠囨倿閿斿墽鐭嗛悗锝堝煐閿燂�???闂佽法鍠曟慨銈吤洪敓�????瀹曟繂鈻庤箛鏇熸闂佺粯鍨归悺鏃堝极閸ヮ剚鐓熼柡鍐ㄦ处椤忕娀鏌￠崱鎰伄缂佽鲸鎹囧畷鎺戭潩閻愵剙�????闂佽法鍠嶇划娆忕暦閹扮増鍊婚柤鎭掑劚閳ь剙娼￠弻銊╁即閻愭祴鍋撻崨濠庢敯闂傚�?�鑳剁划顖炲礉濡ゅ懎纾块柕鍫濐槸绾惧綊鏌涜椤ㄥ棝鎮￠妷鈺傛櫢闁跨噦�????????缂傚倸鍊烽懗鑸靛垔椤撱垹鍨傞柛顐ｆ礀閽冪喐绻涢幋鐐冩艾危閸喍绻嗘い鏍ㄨ壘閹垿鏌熼幓鎺嬪仮婵﹥妞藉畷顐﹀礋閿燂拷?濞呫倝姊虹拠鈥虫灈闁稿﹤鐏濋锝嗙節濮橆儵鈺呮煃閸濆嫸锟???閿熻姤绂嶉悙鐑樷拺缂佸瀵у﹢鎵磼鐎ｎ偄鐏存い顫嫹??
    wire        csr_da;
    wire        csr_pg;
    wire [1:0]  csr_plv;

    //trans_addr to dcache
    wire [31:0] ret_data_paddr;
    wire [31:0] if_pred_addr1;
    wire [31:0] if_pred_addr2;

    wire icache_valid_out;

    wire [18:0] invtlb_vpn;
    wire [9:0]  invtlb_asid;
    wire invtlb;
    wire tlbfill;
    wire tlbwr;
    wire [4:0]invtlb_op;
    wire data_uncache_en;
    wire [31:0]   data_paddr_out;
    wire data_tlb_found_out;
    wire [4:0] data_tlb_index_out;
    wire data_tlb_v_out;
    wire data_tlb_d_out;
    wire [1:0]  data_tlb_mat_out;           
    wire [1:0]  data_tlb_plv_out;
    wire [31:0] tlbehi_out;
    wire [31:0] tlbelo0_out;
    wire [31:0] tlbelo1_out;
    wire [31:0] tlbidx_out;
    wire [ 9:0] asid_out;
    wire [31:0] tlbehi_in;
    wire [31:0] tlbelo0_in;
    wire [31:0] tlbelo1_in;
    wire [31:0] tlbidx_in;
    wire [5:0] ecode_in;
    wire [4:0] rand_index;
    wire inst_tlb_found;
    wire inst_tlb_v;
    wire inst_tlb_d;
    wire [ 1:0] inst_tlb_mat;
    wire [ 1:0] inst_tlb_plv;
    wire [ 9:0] asid_in;

    wire same_page;
    front u_front
    (
    
        .cpu_clk(aclk),
        .cpu_rst(rst),
        .not_same_page(not_same_page),

        .pred_taken(BPU_pred_taken),
        .pi_icache_is_exception1(pi_icache_is_exception1),     
        .pi_icache_is_exception2(pi_icache_is_exception2),
        .pi_icache_exception_cause1(pi_icache_exception_cause1),  
        .pi_icache_exception_cause2(pi_icache_exception_cause2),
        .pc_for_buffer1(icache_pc1),
        .pc_for_buffer2(icache_pc2),
        .pred_addr1_for_buffer(pred_addr1_for_buffer),
        .pred_addr2_for_buffer(pred_addr2_for_buffer),
        .pred_taken_for_buffer(pred_taken_for_buffer),
        .icache_pc_suspend(pc_suspend),
        .inst_for_buffer1(icache_inst1),
        .inst_for_buffer2(icache_inst2),
        .icache_inst_valid1(icache_inst_valid1),
        .icache_inst_valid2(icache_inst_valid2),
        .icache_valid_in(icache_valid_out),

    // *******************
        .fb_flush({flush_o[2],flush_o[0]}), //闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠楅悷鈺侇嚕閸洖鍨傛い鏇炴噹濞堫參姊婚崒姘炬�??閿熶粙宕愰幖浣哥９闁绘垼濮ら崐鍧楁煥閺囩儑锟???閿熺晫绮婚弽顓熺厱妞ゆ劧绲鹃敓锟???缂佸墽鍋擄拷?锟窖呮崲濠靛洨锟??闁稿本绮岄�?�娲煥閻曞倹锟???闂佸憡鍔忛弬鍌涚濠婂牏鍙撻柛銉ｅ妽鐏忛潧顭胯濠線骞忛敓�?????闂佽法鍠曟慨銈吤哄Ο鐓庡灊閿燂�??閸曨偆鍘撮梺纭呮彧闂勫嫰寮查鍕厱闁哄洢鍔屾禍妤呮煛婢舵ê寮慨濠呮缁瑩宕犻埄鍐╂毎闂備焦鎮堕崝�?勬�?�濠靛鍋╅柣鎴ｆ閸楁娊鏌曡箛濞惧亾閾忣偒鍚囧┑锛勫亼閸婃牜鏁繝鍕焼濞达綀顫夐崕鐔封攽閻樺弶澶勯柍閿嬪灴閺屾盯骞橀弶鎴犵シ婵炲瓨绮嶇换鍕閹烘梹瀚氶柤纰卞劮閵徛颁簻妞ゆ挾鍋為崰姗堟�??閿熺瓔鍠曠划娆愪繆濮濆矈妲惧銈嗘⒐濞茬喖骞冨Δ鍛仭闁哄顑欏Λ宀勬⒑閸濄儱校婵炲弶绮撻幊鐐烘焼�?�ュ懐顦х紓浣诡殙濡椼劎鑺辨繝姘拺闂傚牊渚楀Σ鍫曟煕鎼淬�?�鐝柡鍛版硾閳藉顫濇潏鈺嬬床缂傚倸鍊烽悞锕傦�??锟介崶顬＄尨�????閿熻姤锕╁▓浠嬫煟閹邦剚鈻曢柛搴㈡閺岀喖顢欓悾灞惧櫘闂佸湱鎳擄�??锟筋厾绮悢纰辨晬婵炴垼椴搁敍鍫濃攽閻樻鏆滅紒杈ㄦ礋�?�曟垿骞嬮敓�????绾惧湱鎲歌箛鎿冨殫濠电姴鍟伴々鐑芥�?�閿濆簼绨芥い锟??鍔曢—鍐Χ閸℃衼缂備胶濮甸崹鍧�?箖閿熺姵鏅搁柨鐕傛嫹?闂佸搫鐬奸崰鎰焽韫囨稑�?堢憸蹇涘汲閻樼粯鈷戠紓浣股戦幆鍫㈢磼缂佹绠烇拷?锟筋喛顕ч埥澶愬閻橀潧濮堕梻浣告啞閸斞呯磽濮橆兘鏌︽い蹇撴绾捐棄霉閿濆娑у┑鈥虫健閺屾稑螣閻樺弶绁柟鍑ゆ�??闂佽法鍠嶇划娆忕暦閿燂拷?椤㈡瑩宕叉竟顖氭处閻撴洟鏌熼幍铏珔濠碉�??锟藉悑閵囧嫰顢楅�?顒勬偋閹炬剚娼栨繛宸簻缁犱即骞栧ǎ锟??鐏╂い锔规櫆缁绘冻锟???閿熻姤顭囬惌銈吤瑰⿰鍕畺缂佸矉�???????婵犵妲呴崹鐢稿磻閹版澘绠犳繝闈涱儐閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曨敊婵劒绨婚梺鍝勬祩娴滅偟绮旈濮愪簻闁靛骏锟???閿熻棄鎽甸梺璺ㄥ櫐閿燂拷??闂佽法鍣﹂敓�??????闂備椒绱徊鍧楀礂閿燂拷?楠炲啴鍩勯崘鈺佸妳濠碘槅鍨崇划顖炲级閹间焦鈷戦悹鍥ㄥ絻閸よ京绱撳鍛棡缂佸倸绉撮埞鎴�??閿熺瓔浜濇潏鍫濐渻閵堝懐绠伴柣锟??锕崺娑㈠箳濡や胶鍘遍柣蹇曞仜婢т粙骞婇崨顔轰簻闁挎棁鍋愰悾鐢告煛閿燂�??閸犳捇宕版繝鍥х闁绘劖澹嗛惄搴ㄦ⒑缂佹ɑ灏柛濠冪箞�?�寮撮悢铏诡啎闂佺粯鍔﹂崜姘舵偟閺冨牊鈷戞慨鐟版搐閳ь兙鍊濆畷鎶芥晲婢跺﹨鎽曞┑鐐村灦缁姴危閻撳寒娓婚柕鍫濆暙婵″ジ鏌熼搹顐㈠闁告帗甯楃换婵嗩潩閸忓吋娅栨繝鐢靛仦閸ㄨ泛顫濋妸鈺婃晩闁哄洢鍨洪崐鐢告煟閻斿憡绶叉い銉ョ箻閺屾盯鎮╅搹顐ゎ槶闂佸ジ缂氭ご鍝ョ紦娴犲宸濆┑鐘插楠炴姊绘担绛嬫綈鐎规洘锚閳绘柨鈽夐�?鐘插殤濠电偞鍨崹娲偂濞戙垺鏅搁柨鐕傛�??闁诲函缍嗛崜娆撳春锟??鍕叄濞村吋鐟х粔�???鏌＄仦鍓р槈闁宠鍨垮畷鍗炍旀繝浣瑰亝缂傚倸鍊烽悞锕傦�??锟�?�箛娑樼煑闁告劦鐓堝鏍ㄧ箾瀹割喕绨奸柛瀣�??锟介獮鏍垝鐟欏嫷娼戝┑鈽嗗亜閺堫剛鎹㈠☉姘ｅ亾濞戞瑯鐒介柣顓滐�??锟介湁婵犲﹤绨肩花缁樸亜閺囶亞鎮奸柟椋庡Т闇夐悗锝庡亽濞兼棃姊婚敓�????濞佳呮崲閹烘挻鍙忛柣銏℃綄婢跺ň鏀介悗锝庡亞閸樹粙姊虹紒妯忣亪宕㈤弽顓熷殝妞ゅ繐鐗婇悡鏇㈡煛閸屾碍鍋ラ柛娆忓閳ь剝顫夊ú妯兼崲閸儻�????閿熻棄鈽夐姀鈽呮�???????婵犵數濮烽弫鎼佸磻濞戙垺鍋嬮柛鈩冪⊕閸婅埖绻濋棃娑卞剰闁告垹�???閺屾洟宕煎┑鎰﹂梺鍛婂灩婵敻濡甸崟顔剧杸闁规崘娉涢敓�????闂備胶绮幐鎼佸疮閹绢喖绠栫憸鐗堝笒閻愬﹦鎲稿鍥╂／鐟滄棃寮诲☉銏★拷?锟斤�??锟藉壊鍠楁缂傚倷娴囨ご鍝ユ暜閿熺姴绠栭柍杞拌兌閿燂�????缂傚倸鍊搁崐鐑芥嚄閸撲礁鍨濇い鏍ㄧ矋瀹曟煡鏌涢锝囩畼闁哄棴绠撻弫鎾绘晸閿燂�????闂備胶纭堕弲顏嗘崲濠靛棛鏆﹂柟鐑樺灍濡插牊鎱ㄥ鍡楀妞ゅ繐缍婂濠氬磼濮橆兘鍋撻幖浣哥９闁归棿�?佺壕褰掓煙闂傚顦︾痪鎯х秺閺岋綁骞嬮敐鍛呮捇鏌涢妶鍛伃闁哄本鐩獮�???鎳犻澶嬓滈梻浣规偠閸斿秶鎹㈤崘顔嘉﹂柛鏇ㄥ灠閿燂拷?濡炪倖鍔﹂敓�????缂侇噯锟????濠电姰鍨奸崺鏍礉閺嶎厽鍋傛繛鎴欏灪閻撴洟鏌曟径鍫濈仾婵炲懎鎳橀弻娑㈠箻鐠佽櫕鍠氶梺鍝勬湰閻╊垱淇婇崼鏇炲�?�婵☆垳鈷堝Σ褰掓⒒娴ｅ憡鎯堥柡鍫墴閹嫰顢涢悙顏佸亾閿燂拷?瀵挳锟??閳╁啯鐝抽梻浣虹《閸撴繈鎮烽姣硷綁顢楅崒婊咃紳闂佺ǹ鏈悷褔宕濆澶嬬厱闁哄啠鍋撻柣妤冨█婵℃挳宕橀鐓庯拷?锟藉┑鈽嗗灠閻ㄧ兘寮ㄩ搹顐ょ瘈闁汇垽娼у瓭濠电偞娼欓崐鍨嚕椤愩埄鍚嬮柛鈩冪懅椤旀洟姊洪悷閭﹀殶闁稿鍠栭妴鍌炲蓟閵夛妇鍘鹃梺鍓茬厛閸犳寰勯崟顖涙櫢闁跨噦锟???????婵犵妲呴崹鐢稿磻閹扮増鍋傚ù锝堟绾捐棄銆掑顒佹悙闁哄鍠栭弻鐔兼偡閻�?牊鎮欏銈嗘穿缁插墽鎹㈠┑鍡╂僵妞ゆ巻鍋擄拷?锟芥挸妫濆娲箰鎼达絺妲堥柣搴㈠嚬閸ｏ絽顕ｉ崼鏇炲窛濠电姴瀚惁鍫ユ⒑濮瑰洤鐏叉繛浣冲啰鎽ラ梻鍌欒兌鏋柨鏇樺劦楠炲啴宕掗悙鍙夋К濠电偞鍨堕悷銉ф閻愮儤鐓欓梺顓ㄧ畱楠炴劙鏌熼柨瀣仢婵﹨娅ｉ幉鎾礋椤愩垹笑濠电姵顔栭崰鎾诲磹濠靛棭鍤曟い鎰堕檮閻掔》锟???閿熷鍎卞Λ娑㈠储闁秵鈷戦柛婵嗗閺嗗﹪鏌涳�??锟筋偅宕岄柡�?嬬秮閹垽宕ｆ径瀣絽婵＄偑鍊栧ú鈺冨緤閸撗勫床婵犻潧妫鈺傘亜閹捐泛浠掔紒銊ㄥ吹缁辨挻鎷呴崫鍕婵犳鍨垫慨銈夊Φ閺冨牆绠瑰ù锝呮憸閺屟囨煥閻曞倹锟????闂備礁鐤囬～澶愬垂閸ф绠栨繛鍡樻尭缁狙囨煙鐎电ǹ小婵℃鎹囧缁樻媴閽樺鎯為梺闈╃祷閸庨潧鐣疯ぐ鎺戠閿燂拷?閳ь剚绂嶉柆宥嗏拻濞达絽鎲￠崯鐐烘煕閺傝法绠伙�??锟筋喗褰冮埞鎴﹀醇濠靛柊姘舵⒑闁偛鑻晶锟??鏌嶇憴鍕伌闁诡喗鐟╅幊鐘活敆閳ь剟銆傚ú顏呪拺閻犲洩灏欑粻鑼磼鐠囪尙澧曟い鏇秮楠炴牗鎷呴崫銉晪缂傚�?�鍊烽悞锕傦�??锟介崶锟??鍌ㄩ梺锟??绉甸悡鐔煎箹閹碱厼鐏ｇ紒澶屾暬閺屾冻�????閿熺瓔浜濋崳褰掓煟閿濆妫戝ù鐙呯畵閹瑩顢楅�?�???顕ｉ幐搴ｇ瘈闁汇垽娼у瓭闂佺懓鍟跨换锟??銆侀弮鍫熷亹闁汇垻鏁搁敍婊堟煛婢跺﹦澧戦柛鏂跨灱缁參骞掑Δ浣瑰殙闂佹寧绻傞ˇ浼存偂閺囥垻鍙撻柛銉ｅ妽閿燂拷?闁汇埄鍨伴悥濂稿蓟閿涘嫧鍋撻敐鍛暢闁伙絽鐏氶幈銊︾�?閸曨厼绗￠梺鐟板槻閹虫ê鐣烽妸鈺傤棃婵炴垶姘ㄦ婵＄偑鍊戦崹娲偋閻樿尙鏆﹂柛妤冨亹濡插牊淇婇婧炬嫛闁哥偛鐖煎缁樻媴閸濄儳楔濠碘槅鍋勫锟犲箖閻愮儤鏅滈柛鎾楀倻鐟濋梻浣告贡閸庛�?�銆冮崱娑樼厱闁圭儤鍤氳ぐ鎺撴櫜闁告侗鍠栧▓�???姊洪棃鈺佺槣闁告ǹ妫勯悾鐑藉蓟閵夛妇鍘甸梺缁橆殔閻�?﹦娆㈤弻銉﹀仭婵炲棙鐟ч悾鐢告煙椤旂瓔娈滈柡浣瑰姈閹柨鈹戦崼鐔告闂傚�?�绀�?幖顐⑽涳�??锟藉摜涓嶉柟鎹愵嚙缁犳牠鏌ㄩ悤鍌涘?闂佽鍠楅悷鈺佄涢崘銊㈡婵°倐鍋撴い銉﹀哺濮婄粯鎷呴崨濠傛殘闂佽崵鍠嗛崕鎶藉箲閵忋�?�绠涢柡澶庢硶閸樻挳姊虹涵鍛涧闂傚嫬�?�板畷鎴�?箛閻�?牏鍘电紓鍌欑劍閿氬ǎ鍥锋嫹??闂傚倸鍊烽悞锕傛儑瑜版帒鏄ラ柛鏇ㄥ灠閸ㄥ倿姊洪敓�????缁夌敻宕曟惔鈧簻闁哄稁鍋勬禒婊堟煢閸愵亜鏋涢柡�?嬬秮瀵噣宕奸锝庢闂備礁鎼Λ妤咁敄婢舵劖鏅搁柨鐕傛嫹???闂備胶绮�?�鍛涘Δ鍛厺闁圭偓绶為弮鍫濆窛妞ゆ棁顫夛拷?锟藉ジ姊绘担钘夊惞闁哥姵鍔栫粩鐔煎幢濞戞瑦娅栭悗骞垮劚椤︿即鎮￠弴銏℃櫢闁跨噦锟???????婵犵數鍎戠徊钘壝洪妶澶嬫櫇妞ゅ繐鐗嗙粻鏍煕瑜庨〃蹇涘极瀹ュ鐓ユ繝闈涙閿燂拷?閻熸粍鏌ㄩ～蹇曠磼濡偐�????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰�???闂備礁鎼悮顐﹀礉閹存繍鍤曢柟缁㈠枛鎯熼梺闈涚墕濞层劌鈻旈幐搴濈箚闁绘劦浜滈�?顑撅�??锟藉畷鎴�?礋椤撶喎搴婇梺褰掑亰閸犳牕顕ｉ崣澶夌箚闁绘劦浜滈�?顒佹礈閹广垽骞囬懜闈涱伓?闂佽法鍠撻悺�???绂嶉悙鍙傦綁骞囬弶鍧�?敹闂佸搫娲ㄩ崯鍧�?箯濞差亝鈷掗柛灞炬皑婢ф稑銆掑顓ф當閸楅亶鏌涢锝嗙闁绘挻娲熼獮鏍庨敓�????閻忣喗绻涢崣澶嬪唉闁哄备鍓濋幏鍛存偡閺夋娼氶柣搴ゎ潐濞叉牕鐣烽鍕厺閹兼番鍔�?粻锝嗐亜閹捐泛浠︽繛鍛殜濮婂宕掑顑藉亾瀹勬噴褰掑炊閿燂�??绾惧鏌熼悧鍫熺凡闁绘挻娲熼弻娑㈩敃閻樻彃濮庣紓浣插亾闁割偆鍠撶粻楣冩煕閳╁叐鎴犱焊椤撱垺鐓曢柟瀵稿Т鏍＄紓浣虹帛閻╊垶鐛拷?锟筋喗鍊烽柛鎰ㄦ櫅閸濈尨�????閿熺瓔鍠撻崝宥囩矉閹烘柡鍋撻敐搴′簽闁告ɑ鎹囧娲濞戣鲸肖闂佺ǹ瀛╂繛濠囧极瀹ュ拋鍚嬪璺侯儑閸樼敻姊烘导娆戝埌闁兼椿鍨堕崺銏ゅ醇閵夛妇鍘搁梺璺ㄥ櫐閿燂�???闂佸摜濮撮柊锝夊箖妤ｅ啯鏅搁柣妯哄暱娴滈亶姊洪崜鎻掍簼缂佽鍟撮、鏃堝Χ婢跺鎷绘繛杈剧到閹诧繝宕悙鐑樼厽婵°倓绶″▓婊堟煙椤斻劌娲﹂崑鎰舵嫹?閿熻棄澹婇崰鏍�?枔閵娾晜鈷戦柛锔诲弨濡炬悂鏌涢悩鎰佹疁鐎规洘鍔欓幃婊堟嚍閵夈垺�?�介梻浣稿閸嬪棝宕板鍥偨閺夊牄鍔庣粻楣冩⒒閸屾凹鍤熼柣顓熺懄閹便劍绻濋崒銈囧悑閻庤娲樼敮鎺楋綖濠靛鏁勯柦妯侯槷婢规洟姊虹紒妯虹伇濠殿喓鍊濆畷鐢稿礋椤栨稓鍘遍梺瑙勫礃鐏忔瑩宕濆澶嬬厱闊洦姊婚惌鎺楁煛鐏炲墽娲存い銏℃礋閺佹劙宕卞▎妯伙�????闂備礁澹婇崑鍡涘窗閹剧粯鏅搁柨鐕傛嫹?闂傚倸鍊搁崐鎼佹偋婵犲啰鐟规俊銈呮噹绾惧潡鏌熼幍顔碱暭闁绘挻娲熼幃妤呮晲閸涱収鏆㈤梺璺ㄥ櫐閿燂拷??闂傚倷绀�?幖顐ゆ偖椤愶箑绀夐柟瀛樼箥閸ゆ洟鏌熺紒銏犳灍闁稿﹪鏀辩换娑㈠级閹搭厼鍓版繛�?�樼矊婢т粙骞夐幖浣瑰亱闁割偅绻勯悷銊х磼閻愵剙鍔ら柣蹇旂箞閸╃偤骞嬮敂钘変汗闂佸憡鐟ラˇ顖炈囬埡鍛拺缂備焦蓱鐏忎即鏌ｉ埡濠傜仸鐎殿喛顕ч埥澶愬閻樼數鏉搁梻浣哥枃濡椼劎绮堥敓锟???閳ユ牭锟???閿熺瓔鍋嗛敓�????闂佽法鍣﹂敓�?????闂佸憡娲﹂崢浠嬪礆濞戙垺鈷戦柛婵嗗鐎氭壆绱掓径濠勭Ш鐎殿噯锟??????婵＄偑鍊曠换鎰涘☉銏犵疇闁糕剝绋掗埛鎺楁煥閻曞倹锟???濠电偘鍖犻崗鐐☉閳诲酣骞嬮悙�?�橆唶闂備礁�?遍崕銈夛�??锟介幇顔剧闁哄秲鍔庨敓�????闂傚倸鐗婃笟妤呭磿閹扮増鐓涢柛娑卞枤閿燂�??闂佸搫鏈粙鎴﹀煡婢舵劕�???闁绘劕妯婂缁樹繆閻愵亷�????閿熶粙宕曢弻銉﹀殞濡わ絽鍟悡锟??鏌熸潏楣冩�?�闁稿鍔欓弻娑拷?锟介幋婵呯凹濠殿噯绲斤拷?锟芥澘顫忛搹鍦煓婵炲棙鍎抽崜閬嶆⒑閹稿孩纾搁柛銊ョ秺閹�?箖鎮滈懞銉ヤ汗缂傚�?�鐒﹂敋濞存粌缍婇弻锝夋偐閸欏鈹涢梺璺ㄥ櫐閿燂�??????闂傚倸鍊搁崐椋庢濮樿埖鏅搁柨鐕傛嫹??闂傚倷鑳舵灙閻庢稈鏅滅粩鐔煎幢濞嗘劦娼熼梺鍝勫暙閻楀棝宕￠幎鑺ョ厪闊洤锕ラ鍡涙煙妞嬪海甯涚紒缁樼⊕濞煎繘宕滆琚ｆ繝鐢靛仜閹锋垹绱炴担閫涚箚閻庢稒顭囬敓�????闂佹悶鍎崝搴ㄥ储闁�?秵鈷戦悷娆忓閸斻�?�銇勯弴銊ュ箻缂侇喖顭烽幃娆撴�?�濡厧骞嶆俊鐐拷?锟藉褰掑磿閹惰棄鍌ㄩ柟缁㈠枟閻撴稑霉閿濆毥褰掑汲閿濆鏅搁柨鐕傛嫹??濠碉紕鍋戦崐鏍暜閹烘柡鍋撳鐓庡籍鐎规洘鍨块崺锟犲川椤�?儳骞楅梻浣侯攰閹活亞寰婃ィ鍏寰勯幇顓犲弮闂佸憡鍔︽禍婊堝几濞戙垺鐓涢悘鐐靛亾�???鍐挎�??閿熻姤婢橈拷?锟筋剟鍩ユ径濠庢建闁糕剝锚閺嬬娀姊婚崒娆戭槮闁硅绻濋垾锕傚炊閿燂拷?閺嬩線鎮归崶褎鈻曟繛鍏肩墬缁绘稑顔忛鑽ょ泿闂佸湱顢婇崺鏍Φ閸曨垰绠婚悗鐢电《婵洭鏌ｆ惔銏㈩暡闁烩晩鍨伴～蹇撁洪鍕獩婵犵數鍋炵敮鈺傜椤忓懍绻嗛柛顐ｆ�?缁犵懓霉閿濆懏鎲搁柣锝呮惈閳规垿顢欐慨鎰捕闂佺ǹ顑嗛幑鍥�?蓟閳╁啯濯撮悷娆忓绾炬娊姊虹拠鈥虫�?闁哄懐濮撮悾宄拔熸總钘夋贡閳ь剨缍嗘禍娆愮珶閺囥垺鈷戦柛鎾瑰皺閸樻盯鏌涳拷?锟筋亝鍤囷拷?锟芥洩锟??缁犳盯寮崜褏鐣炬俊鐐�??锟介悧妤冨垝閿燂�??閺侇喚鎹勬總鐣屾�?楗即宕奸姀銏℃瘒闂備浇顕栭崰妤咃拷?锟介崨杈剧稏婵犻潧顑嗛崐鐑芥煥閻曞�?�锟???闂佽法鍣﹂敓�??????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠掗弲鐘荤嵁閹捐绠抽柡鍐╁灥閺咁亪姊婚崒姘炬�??閿熶粙宕愰幖浣哥９濡炲娴烽惌鍡椕归敐鍫燁仩閿燂�??婵犲倵鏀介柣妯垮紦鏉╄绻涢幋娆忕仼闂佽￥鍊濋弫鎾绘晸閿燂拷??????闂傚倸鍊烽悞锔兼�??閿熺獤鍏犲搫顓兼径濠勶紱闂佺懓澧界划顖炴偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺戞倯闁靛洤瀚伴弫鎾绘晸閿燂�???缂傚倸绉撮敃顏勵嚕閿燂拷????闂佽鍑界紞鍡涘礈濞戙垺鍎婇柛顐犲劜閸婄敻鎮峰▎蹇擃仾閿燂拷?閳ь剟鎮楃憴鍕�?闁告挾鍠栧畷娲Ψ閿燂拷?缁剁偛鈹戦悙顏勭仾婵﹤缍婇獮蹇涘川閺夋垵绐涙繝鐢靛Т鐎氼亝绔熼弴鐐╂�?闁绘ê鐏氶弳鈺佲攽椤旂偓鏆い銏＄懇�?�粙顢�?悙鐢靛炊闂備礁鎼粙�???宕㈡禒�?�柧婵犻潧顑嗛悡蹇撯攽閻愯尙浠㈤柛�???顨婇弻鈽呮嫹?閿熺瓔浜炴晥闂佸搫琚崝�?勫煘閹达箑骞㈡俊顖欒濡茶鲸淇婇悙顏庢嫹?閿熶粙宕戦崨顒兼椽鎮㈤悡搴ゆ憰闂佺粯鏌ㄩ崥�?�磹缂佹ü绻嗘い鏍ㄧ矊閸斿銇勯敓锟???濞茬喎顫忛搹鍦＜婵☆垵宕甸崣鍡涙⒑閸涘﹨澹樻い鎴濐槸閻ｇ兘鎮界粙璺唺濠德帮拷?锟介懗鍫曞储椤忓牊鈷戦柛鎾村絻娴滄繄绱掔拠璇ф�??閿熶粙銆佸Δ鍛潊闁靛骏锟???閿熸垝绮￠梻浣瑰缁诲�?�藝娴兼潙鐓曢柟鐑橆殕閻撴洟鎮橀悙鏉戠濠㈣锕㈤弻宥堫檨闁告挻鐩畷锟??顫滈�?顒勭嵁婵犲伣鏃堝川椤斿吋鐤傞梻浣圭湽閸ㄥ綊宕ラ埀顒傜磼椤旇姤灏︽慨濠傤煼瀹曟帒鈻庨幋婵嗩瀴闂佽娴烽悷鎶藉礂閻樿崵绱扮紒鐘崇☉閳藉螣绾拌鲸�???闂備礁鎲″ú锕傚礈濞嗘劗顩峰┑鍌氭啞閳锋垹绱撴担濮戭亪鎮橀崡鐐╂斀妞ゆ柨鎼埀顒佺箓閻ｇ兘骞嬮敓锟???鎯熼梺鍐叉惈閸婄敻骞忔繝姘拺闁告挻褰冩禍鐐烘煕閻樿櫕宕岄柛鈹垮劜�?�板嫰骞囬鐘插箺闂傚⿴鍋勫ú锕傚箹椤愶妇鍙曟い鎺嶇劍閸欏繐鈹戦悩鎻掓殲闁靛洦绻勯�?顒冾潐濞叉鍒掗幘鑽ゅ祦闁规崘顕х粻绛规嫹?閿熷鍎卞ú锕傚疾婵傚憡鈷掗柛灞剧懅椤︼箓鏌熼懞銉х煁闁逛究鍔戝鍫曞箠閵娧勫殌闁伙綇绻濋獮宥夋惞椤愩�?�鍋撴繝姘拺闂傚牊绋撶粻鐐烘煕婵犲啰澧碉拷?锟芥洘鍔栫换婵嗩潩椤撶姴骞堥梻锟??娼ч敓�????缂佽尪濮ゆ穱濠囧礂缁楄桨�??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕敐鍡╂綉闂佸搫妫旈崡鍐差潖缂佹ɑ濯撮柛娑㈡涧缂嶅﹪銆侀弽顓炲�?�婵炴垶顭囬澶愭⒑閹肩偛鍔撮柛鎾寸懇閹锋垿鎮ら崒娑橆伓?闂佽法鍠庨～鏇㈠磿闁�?秵鍋嬫繝濠傚枤閻庡爼鏌曟繛鐐珕闁抽攱鍨块弻娑樷槈濮�?牊鏁鹃柣蹇撶箣閸楁娊寮婚敐澶嬪亜闁哄鍨甸～鍥煥閻曞�?�锟???????婵＄偑鍊曠换鎰矓閻㈢鍋撻棃娑氱劯婵﹥妞藉Λ鍐ㄢ槈濮橆剦鏆繝纰樻閸嬪懐绮欓幒锟??鐤鹃柛顐ｆ礃閻掔》锟???閿熷鍎卞Λ娑㈠储閿燂�?????闂佽法鍣﹂敓�??????濠电偛顕敓�????濞存粌鐖煎濠氭偄绾拌鲸鏅╅梺绋跨箰椤︻垱绂嶆ィ鍐╃厸闁稿本锚閸�?粍銇勯銏⑿㈤柍瑙勫灴椤㈡瑧绮碉�??锟筋偆鏆ユ繝纰樻閸嬪懘鎯勯姘辨殾妞ゆ帒�?�崑銊╂煕濞戞﹫鍔熼柛妯圭矙濮婅櫣绱掑鍡欏姺闂佺ǹ绨洪崐婵囦繆閹绢喖绀冩い鏃囨娴�?垶姊洪柅鐐茶嫰婢ф挳鏌℃担绋挎殻鐎规洘甯掗～婵嬪箟鐎ｎ剙鎯炴繝鐢靛Х閺佹悂宕戦悙鍝勫瀭妞ゆ牜鍋涢崹鍌涚箾瀹割喕绨奸柛瀣�??锟介弻锟犲炊閵夈儳浠肩紓浣哄Т缂嶅﹪骞冮敓�????閳藉鈻庡Ο鐓庡Ш闂備礁鐤囧Λ鍕囬悽鍛婃櫢闁跨噦�??????缂傚倷绶￠崰鏍儗娴ｅ浜瑰〒姘ｅ亾婵﹥妞介獮鏍倷閹绘帒螚闁诲骸绠嶉崕閬嶆偋閸℃稑绠氶柛顐ゅ枍缁诲棝鏌曢崼婵囨悙閸熸悂姊虹粙娆惧剳闁稿鍊濋悰锟??骞嬮敓锟???閻愬﹥銇勯幒鎴�??閿熺晫绮婇敃鍌涒拺闁革富鍘奸崝�?�亜閵娿儲鍣介柣姘劤椤撳吋寰勶拷?锟筋剙骞堥梺璺ㄥ櫐閿燂拷??????闂傚倷绀�?幉鈥愁潖瑜版帒鍨傞柣銏ゆ交缂嶆牠鐓崶銊р姇闁诡垳鍋ら幃宄扳枎韫囨搩浠奸梺缁樼箑閸�?啿顫忓ú顏咃拷?锟介柦妯侯槸婵倕鈹戦悙鍙夊櫤婵炶尙鍠栭獮鍐ㄎ熸笟顖氭�?�闂佸憡绮堥悞锔兼嫹?閿熻棄鐭傚娲濞戞艾顣洪梺鍝ュ櫏閸嬪懏绌辨繝鍐檮闁告稑锕﹂崢鐢告⒑閹勭闁稿鎹囬幊鎾诲锤濡や胶鍘告繛杈剧悼閹虫挻鎱ㄥ澶嬬厵妞ゆ梻鏅幊鍐婢舵劖鏅搁柨鐕傛�?????闂傚倸鍊峰ù鍥敋瑜斿畷娆撴偩鐏炵晫绛忔繛瀵稿Т椤戝棝宕愰懜鍨弿婵☆垱瀵х涵楣冩煟閵堝鐣洪柡灞炬礉缁犳冻锟???閿燂�??锟藉煐閿燂拷??闂佽法鍠嶇划娆撳春濞戙垹绠ｉ柣妯兼暩閿涙粓鏌ｆ惔顖滅У闁稿�?�伴弫鎾绘晸閿燂�?????闂備浇顫夐鏍窗濮樺崬顥氬┑鍌氭啞閻撳繐鈹戦悙鎻掔殹闁瑰嚖�????闂佽法鍠嶇划娆撳箚鐏炶В鏋庨煫鍥э攻閿燂�??闂備焦鏋奸弲娑㈠疮椤栫偛纾归柟鎵閻撴洟鏌嶉崫鍕靛剳缂佲檧鍋撻柣搴ゎ潐濞叉鏁�?幒鏇犱簷濠电偠鎻徊鑺ョ珶婵犲啫顕遍柡宥庡幗閳锋帡鏌涚仦鍓у暡闁瑰嚖锟???闂佽法鍠撻弲顐ゅ垝閸儲鏅搁柨鐕傛嫹?濡ょ姷鍋涢ˇ鐢稿极瀹ュ绀嬫い鎺嗗亾閹兼潙锕铏圭矙閹稿孩鎷辨繝銏ｎ潐濞茬喎鐣烽幋锟??绠婚柟棰佺劍閸嶇敻姊虹紒妯诲碍婵炴挳�?辩粋鎺楀箹娴ｅ厜鎷洪梺鍦�?瑰ù椋庣不閿燂�??閺屾冻锟???閿熷鍔岄埀顒佺箓椤曪綁顢曢敓锟???�???鍐┿亜閺冨洤浜归柨娑欑矊閳规垿鎮欓弶鎴犱桓闂佺厧缍婄粻鏍偘閿燂�??瀹曞ジ濡烽敂瑙勫濠电偠鎻敓锟???濠殿喓鍊�?☉鐢稿醇閺囩喓鍘遍梺鎸庣箓缁绘帡鎮鹃崹顐闁绘劘灏欑粻濠氭煥閻曞�?�锟??????闂傚倸鍊搁崐鎼佸磹閻戣姤鍊块柨鏇烇拷?锟界粻鏍煕椤愶絾锟??閿燂�??婢舵劖鍊堕柣鎰暩閹藉�?�鏌ｉ幒宥囩煓闁哄被鍔戦幃銏ゅ传閸曟埊缍�?弻娑虫嫹?閿熺瓔鍊栭幋�???桅闁告洦鍨伴崡鎶芥煥閻曞倹锟???婵炲瓨绮撶粻鏍箖濡ゅ啯鍠嗛柛鏇ㄥ墰椤︺劑姊洪幐搴㈢８闁搞劋绮欐俊�?�樻媴缁洘鐎婚梺鐟扮摠缁诲啴鎮楅幎鑺ョ厸濠㈣泛锕︽晶鎴︽煕閺傛寧鎹ｇ紒顔芥閺屽棗顓奸崱蹇斿闂備胶枪閺堫剟鎮疯缁綁寮�?�?顒傛崲濞戞瑦濯撮柛鎰�?级婢跺嫰鏌涳�??锟筋亶鍎旈柡灞剧洴閸╁嫰宕橀浣诡潔缂傚倷鑳舵慨閿嬬箾閳ь剟鏌￠敓�????閸犳牕顕ｉ崼鏇炲瀭妞ゆ棁鍋愶�??锟藉ジ姊绘担瑙勫仩闁稿海鍎ょ粋宥囨崉娴ｆ洜鍠栧畷鐔碱敃閻斿憡鏉告俊鐐拷?锟藉濠氬Υ鐎ｎ�?�娑橆潩椤撶姷顔曢梺鍛婄矊閸熶即骞冩總鍛婄厱闁圭儤鎸哥粭鎺楁煃鐠囨煡鍙勬鐐差儔閹瑩鎳犻濠勭闂傚�?�鍊风欢姘焽瑜戦崳褰掓煟韫囨洖浠╁┑顔猴拷?锟藉鎶筋敍閻愮补鎷婚梺绋挎湰閻旑剟骞忛敓锟????闂佽法鍠撻弲顐ゅ垝閸儲鏅搁柨鐕傛嫹?濡ょ姷鍋涢ˇ鐢稿极閿燂�??????闂傚倷鑳剁涵鍫曞礈濠靛牏鐭欓柟�?�稿Х閻棝鏌涢幇闈涙灍闁绘挶鍎茬换婵嬫濞戞瑯妫″銈冨劤閿燂拷?闁哄矉锟?????闂備礁婀遍埛鍫ュ磻婵犲洤鏄ラ柣鎰惈缁狅綁鏌ㄩ弮鍥棄濞存粌�?辩槐鎾诲磼濞嗘垵濡介柦鍐憾濮婂搫鈻庨幆褍绠瑰銈庝簻閸熷瓨淇婇崼鏇炲�?�婵°倕鍟╁ǎ顔界節绾版ɑ顫婇柛�?�噽閹广垽宕煎┑鍫熸闂佸憡绻傦拷?锟窖兾ｉ崼銉︾厪闊洦娲栧暩濡炪倖鏌ㄩ敃顏勵潖濞差亜鎹舵い鎾跺仒缂傛捇姊洪崨濠冪叆闁活剝鍋愬Σ鎰版倷鐎靛摜鐦堥梺鎼炲劀閸曨厸鍋撻鍕拺闁革富鍘奸。鍏肩節閵忊槄鑰块柡灞筋儔�?�曞爼顢楁担鍝勫箺闂備礁鎼ú锔惧枈�?�ュ＆鍥�?�閼恒儳鍘卞┑鐘绘涧濞村倸鈻撳⿰鍕弿濠电姴鍊归幆鍫ュ极閸儲鐓曢柕澶嬪灥閹冲孩鎱ㄩ崼鏇熲拻濞达�?顫夐崑鐘绘煕閿燂�??閸ㄥ墎绮嬪澶婇唶闁哄洨鍋熼悾楣冩⒑閸涘﹥澶勯柛銊ャ偢�?�偄顓兼径瀣幗闂佸綊鍋婇崹浼存嫊婵傚憡鐓欓柤鎭掑劜锟??瀣叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚�?�鑳剁划顖烇�??锟介崨顖�?亾濮樼厧骞樼紒顔碱儏椤撳ジ宕煎☉妤佺潖闂備礁�?遍崕銈夊箰妤ｅ啫鍌ㄩ柣銏犳啞閳锋垹绱撴担濮戭亪鎮�?敃鍌涘珔闂侇剙绉甸悡鍐⒑閸噮鍎忔繛鎼櫍閺岋�??锟界暆鐎ｎ剛鐦堥悗瑙勬礋娴滃爼宕洪埄鍐╁鐎瑰嫮澧楅悗鍐测攽閻樻剚鍟忛柛鐘崇墵閺佸啴濡搁妷銏★拷?锟介梺鎸庣箓椤︻垳绮婚鐐寸厽婵☆垱顑欓崵娆撴煟韫囨柨鈻曢柡灞熷棛锟??闁挎繂鎳嶇花鑺ョ箾鐎涙鐭庨柛鈺傜墱閹广垹鈹戦崼婵囷�??锟芥繝銏ｆ硾閻ジ鏁嶉悢鍏尖拺缂佸顑欓崕鎰亜椤撶偞鍠橈拷?锟芥洘宀搁獮鎺楀箣閿燂拷?閻庡姊虹憴鍕姢闁哥喎娼￠幃妤咁敇閻斿墎绠氶梺闈涚墕缁绘帡宕氭导�?�樼厱闁绘洑�?�?悘锔兼嫹?閿熺瓔鍠楄ぐ鍐煘閹寸姭鍋撻敐搴′簽闁告﹢浜堕弻锝堢�?閺囩偘鎴烽梺绋款儐閹瑰洭骞嗛崘顔肩闁绘劦浜欑花濠氭⒑閸濆嫸�????閿熺晫浜搁崨瀵稿彆妞ゆ帊鐒﹂崣蹇撯攽閻樻彃鏆為柕鍥ㄧ箘閳ь剝顫夊ú婊堝礂閿燂�??閵嗕礁顫滈埀顒勫箖濞嗘挸绾ф繛鍡欏亾椤ワ繝姊婚崒姘炬嫹?閿熺晫绮堥敓�????楠炲鏁撻悩鑼唶闁荤姴娲╃亸娆撳汲閸℃稒鐓欓梻鍌氼嚟椤︼箓鏌★�??锟解晝绐旈柡�???鍠栧畷婊嗩槾閻㈩垱鐩弻锟犲川椤�?枻锟???閿熶粙鏌＄仦璇插闁诡喓鍊濆畷鎺戔槈濮楀棔锟????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠掗弲鐘荤嵁閹捐绠抽柡鍐╁灥閺咁亪姊婚崒姘炬�??閿熶粙宕愰幖浣哥９濡炲娴烽惌鍡椕归敐鍫燁仩閿燂�??婵犲倵鏀介柣妯垮紦鏉╄绻涢幋娆忕仼闂佽￥鍊濋弫鎾绘晸閿燂拷??????闂傚倸鍊烽悞锔兼�??閿熺獤鍏犲搫顓兼径濠勶紱闂佺懓澧界划顖炴偂閸愵喗鐓㈡俊顖欒濡牊淇婇幓鎺戞倯闁靛洤瀚伴弫鎾绘晸閿燂�???缂傚倸绉撮敃顏勵嚕閿燂拷????闂佽鍑界紞鍡涘礈濞戙垺鏅柣鏂垮悑閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曞礈瑜忕壕鏂ゆ嫹?閿熷鍎遍幊蹇浰夐悙鐢电＜闁稿本姘ㄦ晥闂佽鍠楃划鎾诲箰婵犲啫绶為敓�????婵犲倹鏆╅梻鍌氾�??锟藉ù鍥�?枖閺囥垺鏅搁柨鐕傛嫹????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏ⅵ闁稿﹥顨堢划娆掔疀濞戞瑯妫呭銈嗗姂閸ㄧ儤寰勯崟顖涚厵鐎瑰嫰鍋婇崕蹇涙偂閵堝棎浜滈煫鍥ㄦ尵鏍￠梺鍝勬噺缁挸顫忓ú顏勫窛濠电姴鍟ˇ鈺呮⒑閸涘﹥灏伴柣鐔濆懎鍨濆┑鐘叉处閸ゅ鏌涜箛鎾存喐缂佺姵宀稿铏圭磼濡搫袝婵炲瓨绮嶇划鎾诲春閳ь剚銇勯幒宥堝厡濠⒀冪仛椤ㄣ儵鎮欓弶鎴濐潔闂�?潧鐗炵紞浣哥暦閿燂拷?婵℃瓕顧傜紒杈哺缁绘繈鎮介棃娑楁勃闂佹悶鍔岄悥濂稿箖閻戣棄围闁搞儯鍔屾惔濠囨⒑缁洖澧叉い顓炴川缁骞橀崨顔碱伓?闂佽法鍠曞Λ鍕珶婵犲洤绐楅柡鍥╁Ь婵啿鈹戦崒姘暈闁绘挸鍟村娲垂椤曞懎鍓伴梺璇茬箲閹告娊寮婚敓鐘虫櫢闁跨噦锟???闂佸摜濮甸悧鐘荤嵁婵犲洤�???妞ゆ挾鍋熼崢鍛婄箾鏉堝墽绉い銉︽崌楠炴垿寮撮悙鈺傛杸闂佺粯蓱椤�?牠寮抽鐐寸厓鐟滄粓宕滃┑鍡忔�?�闁哄洢鍨圭壕濠氭煏婢跺棙娅嗛柣鎾寸洴閹﹢鎮欓惂鏄忣潐閺呭爼寮婚妷锔惧幍閻庣懓瀚晶妤呭闯娴犲鐓欓柛娆忣槹鐏忥讣�????閿熻姤娲滈崰鏍�??锟介弴銏″亜闁炬艾鍊搁ˉ姘舵⒒娴ｇ瓔娼愬鐟版閺呰泛螖閸涱喖�???????闂備礁鎼ú銊╁磻閻愬搫绠归柟閭﹀劒瑜版帗鍋戦柛娑樼摠椤庡秶绱撴担铏瑰笡闁烩晩鍨堕獮鍐焺閸愨晛鍔呴梺鎸庣箓濞村�?�宕拷?锟筋亖鏀介柣妯活問閺嗩垶鏌涢幘�?�哥疄闁诡喗妞藉鎾煑閸濆嫭鍠樻鐐达耿椤㈡瑩鎮剧仦钘夌闂傚倷鐒︼拷?锟窖兠哄澶婄；闁瑰墽绮悡鐔兼煥閻曞�?�锟???濠碘槅鍋呯换鍫濈暦濞差亝鍊烽柛婵嗗椤撴椽姊洪幐搴⑩拻缂侇噮鍨跺鏌ュ煛閸涱喒鎷洪梺鍛婄箓鐎氭悂骞忛敓锟????????缂傚倸鍊风粈浣规櫠鎼淬劌鏋侀悹鍥ф▕濞兼牗绻涘顔荤盎鐎瑰憡绻傞埞鎴︽偐閼碱剛�????闁荤姵浜介崝搴ｅ婵傚憡鐓熸俊顖濇閿涘秴顭胯娴滎亪寮婚敐澶嬫櫜闁搞儜鍐ㄧ�???闂傚倷绶氬褔鎮ч崱妞㈡稑螖娴ｄ警娴勫┑鐐叉▕娴滄繈鍩涢幋锔界厱婵炴垶锕崝鐔兼煃閽樺锟??闁硅櫕绻傞悾婵嬪礋椤掑�?�骞嶉梻浣圭湽閸娿�?�宕归柆宥庢晜闁绘鏁哥壕濂稿级閸稑濡斤拷?锟芥洖鐬奸埀顒冾潐濞叉鏁幒锟??鐓濋幖娣�?妼缁狅絾绻濋棃娑欙紞闁诲孩鎸冲濠氬磼濞嗘垵濡介柣搴ｇ懗閸愵亝娈曢梺褰掓？锟??�???鎷戦悢鍏肩叆婵犻潧妫涙晶銏ゆ煥閻曞�?�锟???闂傚倷娴囬～澶愬磿閹惰姤鍋柛銉墮閺勩儵鏌ｉ幇顔煎妺闁抽攱鍨块幃妤呭捶椤撶儑锟???閿熻姤绻涢崗鐓庡闁哄本鐩俊鎼佸Ψ閿燂拷?娴犳挳姊洪棃娑欘棛閿燂拷?閿燂�??閸┿垺鎯旈妸銉ь啋闂佸搫顦伴崹宕囧垝閿熺姵鈷戦悹鍥ㄥ絻椤掋垻绱掞拷?锟筋偄娴�?柡浣割儔閺佹捇鏁撻敓�????????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏缂佹煡绠栧鏌ヮ敂閸啿鎷洪梺鍦瑰ù椋庣不閹炬番浜滈柨鏃囨硶閻瑱�????閿熺瓔鍣�?崑濠傜暦閿燂�??椤㈡瑩鎮剧仦钘夋辈闂傚�?�绀�?幖顐�?疮椤愶箑纾归柣鐔稿閺嬪秹鏌￠崶銉ョ仾闁绘挻娲熼弻锟犲磼濠靛洨銆婇梺绯曟櫔缂嶄線寮婚悢纰辨晩缂佹稑顑嗛悿�???姊虹紒妯圭繁闁革綇绲介悾鐤亹閹烘繃鏅╅梺缁樻尭鐎垫帒顭囧☉妯锋�?闁绘ɑ顔栭弳顖涗繆閹绘帗鍤囷拷?锟芥洘鍨垮畷顭掓�??閿熻姤锚娴狀參姊洪棃娑辨Т闁哄懏鐩幃鈥斥攽閹炬潙�????闂佽法鍠庨～鏇㈠磿闁�?单鍥敍閻戝洨绋忛梺鍛婄☉閻°劑鎮¤箛娑欑厱妞ゆ劧绲跨粻鏍ㄣ亜閵夛箑鐏撮柡锟??鍠栭弻顭掓嫹?閿熺瓔鍋佹禒銏ゆ⒑閸濆嫮鐒跨紓宥勭窔楠炲啴鍩￠崨顓狀槯闂佸憡绋掑锟??鎮炴繝姘拻濞达絽鎲￠崯鐐烘煛鐏炶濮傞柟宕囧枛椤㈡盯鎮欓懠�???骞掗柣搴＄畭閸庨亶藝椤栨粎涓嶆繛鎴欏灪閻撶喖鏌ㄩ悤鍌涘?闂佺粯顨呯换妯虹暦閵忋�?�鍋ㄩ柛娑樑堥幏娲⒑閸涘﹦鈽夐柨鏇橈拷?锟介幃锟??鎮㈤崗鑲╁幈婵犵數濮撮崯鐗堟櫠闁�?秵鐓冪憸婊堝礈濮樿埖鏅搁柨鐕傛嫹????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙宸富闁靛牆妫楃粭鎺楁煥閺囶亜顩紒顔界懆缁犳盯寮崒婊呮闂備線娼ф蹇曞緤閸撗勫厹闁绘劦鍏欐禍婊堟煙鐎涙绠栭柛鐘筹�?�閺�?喖顢欓悙顒佹瘓閻庤娲栭妶绋款嚕閹绢喗鍋勯柛婵嗗缁犵偤姊婚崒娆戝妽闁哄銈稿鎻掆槈閵忕姷鐓戦梺鍦濠㈡绮婚敐鍡欑瘈闂傚牊绋戦弳鐐烘煟鎼淬垺銇濇慨濠呮缁辨帒螣韫囷絼閭�??锟芥洏鍨藉浠嬵敃閿濆懎绨ラ梻浣虹�?�閸撴繄绮欓幒妤佸亗闊洦绋掗悡鏇熴亜閹板墎鎮肩紒鐘崇墵閺屾盯鏁愰崱妯镐虎闂佸搫鏈惄顖炲极閹版澘骞㈡俊顖炴櫜閾忓酣姊绘担鍛婃儓闁哄牜鍓涚划娆撳箻鐠囪尙鍔﹀銈嗗笒閿曪妇绮旈棃娴㈢懓饪伴崟顓犵厜闂佽法鍣﹂敓锟??????婵犵數鍋熼妴瀣箯閿燂拷??闂佽法鍠撻悺鏃堝吹閺囩偐�?介柣妯虹枃婢规﹢鏌涘Δ浣糕枙闁哄矉缍佸锟??宕奸锝庢缂傚倷鐒﹂崝妤呭磻閵堝拋娼栭柧蹇曟嚀鐎垫煡鏌￠崶鈺佷粶闁冲嘲顦甸弻锕傚礃椤旂粯鍠氶梺鍝勭焿缁蹭粙鍩為幋锟??鐐婇柕濞у本效濠电姵顔栭崰鏍晝閵娿儮鏋嶉柨婵嗘处椤洟鏌熼悜妯烘闁绘梻鍎わ�??锟芥岸鏌涘▎蹇ｆЧ妞ゆ柨鍊垮濠氬磼濞嗘埈妲梺纭呭Г缁秹骞堥妸鈺傚仺闁告稑锕ゆ禍閬嶆⒑缂佹◤顏勎熸繝鍥у惞闁哄洨鍋愰弨浠嬫煟濡櫣锛嶆い锝嗙叀閺岋繝宕ㄩ鏂ゆ�??閿熶粙鏌″畝瀣埌閾伙綁鏌涢…鎴濇灓婵絻鍨藉娲箰鎼达絺濮囩紓渚囧枛閻倿宕洪悙鍝勭闁挎棁妫勯�?顒傚厴閺屸剝寰勶�??锟筋亞浠兼繛瀵稿У閹倸顫忓ú顏勭閹兼番鍨婚敍鏇㈡⒑閸濆嫭鍣藉┑顔芥尦閹箖鎮滈懞銉ヤ缓缂佸墽澧楅敋濞存粓绠栭弻銊モ攽閸℃冻锟???閿熶粙鏌★拷?锟筋剙鏋涢柡灞界Ч閺岊煉锟???閿熺瓔浜炴导�?勬⒑閸濆嫭婀扮紒瀣灴閸╃偤骞嬮敓锟???�???瀣亜閹扳晛鐏╂い顐ｆ崌濮婄粯鎷呴崨濠冨創濡炪�?�鍨靛Λ妤勭亱闂佸憡鍔﹂崰鏍嫅閻斿摜绠鹃柟�?�稿仜閻掑綊鏌涳�??锟筋偅宕岄柡浣瑰姍�?�曟﹢濡搁妷顕嗘�??閿熶粙姊婚敓�????閳ь剛鍋涢懟顖涙櫠椤栨粎纾奸悹鍥ㄥ絻閳ь剙娼￠妴浣割潩閼稿灚娅滈梺绯曞墲閻熝囨儊閸績鏀芥い�???鏋绘笟娑㈡煕濡寧顥夐柍璇茬Т楗即宕奸悢鍙夊闂備礁鎲￠幐鏄忋亹閸愨晝顩查柡宥庡幗閻撴洟鏌曟繛鍨姶闁绘捁鍋愰埀顒侇問閸犳牠鎮ユ總鍝ュ祦闁哄秲鍔嶆刊鎾煕韫囨搩妲归悗姘偢濮婄粯鎷呴崨濠呯闁哄浜濈换娑㈠箻椤曞懏顥栫紓渚囧枛椤兘鐛Ο鑲╃＜婵☆垳鍘ч獮宥夋⒒娴ｅ憡鍟為柛锟??顭囨禍绋库枎閹寸姳绗夋繝鐢靛У绾板秹鎮￠敓�??????婵犵數鍋�?崠鐘诲炊瑜忛崢鎾⒑閻熼偊鍤熷┑顕呭弮�?�曟垿骞樼紒妯绘珳闁硅偐琛ラ�?顒冨皺閻栭亶姊绘担鍝ョШ閿燂拷?閸楃儐娓婚柦妯侯樈濞兼牗绻涘顔荤盎鐎瑰憡绻傞埞鎴︽偐閹绘帩�???闂佷紮绲块弫濠氬蓟閿濆棙鍎熼柕蹇曞Т濮ｅ牓姊洪棃鈺冪Ф缂傚秳绶氶弫鎾绘晸閿燂�?????闂備礁鎼懟顖毼涘Δ鍜佹晣濠靛倻枪楠炪垺绻涢崱妤冪缂佺姷鍋ゅ濠氬磼濞嗘帒鍘＄紓渚囧櫘閸ㄧ敻骞楅锔解拺缂備焦蓱閹牏绱掔紒妯肩畵闁伙絿鍏橀弫鎰緞婵犲嫷妲规俊鐐�??锟介悧妤冪矙閹捐鍌ㄩ梻鍫熶緱濞撳鏌曢崼婵囶棡缁惧墽鏁婚弻娑虫�??閿熺瓔鍋呯亸鐢电磼鏉堛劌娴柟顔规櫅閻ｇ兘宕惰閹蜂即鏌ｆ惔銏╁晱闁革綆鍣ｅ畷鎴炵節閸モ晛绁�?┑鈽嗗灥閸嬫劗澹曢崗闂寸箚妞ゆ牗绻冮妴鍐╂叏鐟欏嫷娈滄慨濠勭帛閹峰懘鎸婃径澶嬬潖闂備礁鍟块崲鏌ユ偋閹惧磭鏆︽繝濠傜墛閸嬪嫰鏌涜箛鏇炲付濞寸姵甯�?�娲偡閺夊簱鎸冪紓渚囧櫘閸ㄥ爼宕哄☉銏犵闁圭偨鍔岀紞濠囧极閹版澘宸濇い鏂垮悑濞堟﹢姊洪懡銈呅ｉ柛鏂炲懏宕叉繝闈涙－閸ゆ洟鏌熼梻瀵歌窗闁轰礁鍊块弻娑㈠灳瀹曞洨顔囨繛瀛樼矒缁犳牠寮诲☉銏℃櫆閻犲洦褰冪粻濠氭⒑闂堟稒顥滈柨鏇ㄤ邯瀵鏁撻悩鎻掔獩濡炪�?�鐗楅崺鍐几閸涘瓨鍊甸悷娆忓�???鍐╀繆閻愭壆鐭欙�??锟筋噮鍋婇獮妯肩磼濡桨姹楅梻浣藉亹閳峰牓宕滈妸褎顫曢柛娆忣槺閿燂拷?闂佹眹鍨藉褍鐡梻浣瑰濞插繘宕愬┑�?�祦闊洢鍎查敓锟????闂佽法鍠撻悺鏃堝窗閺嶎厽鍋い鏇�?亾妤犵偞鐗曡彁妞ゆ巻鍋撳┑鈥茬矙閺屽秹鏌拷?锟筋亞鐟ㄩ梻鍥ь樀閺屻劌鈹戦崱妯烘闂佸摜鍠撻崑銈夊蓟閻旂⒈鏁嶆慨妯哄船閿燂拷?闂備線娼уú銈忔�??閿熸垝鍗冲顐﹀磼閻愭彃鐎銈嗘閸嬫劙濡堕敓�????閺岋絾鎯旈妶搴㈢秷濠电偛寮堕悧婊呮閻愬锟??闁搞儜鍛毇闂備椒绱徊浠嬫儔婵傚憡鍎楁繛鍡樻尰閸嬶綁鏌熼鐔风瑨濠碉拷?锟芥健閺岋繝宕遍埡浣峰枈濠殿喖锕︾划顖炲箯閸涘瓨鍊绘俊顖滃劋閻ｎ剚淇婇悙顏庢�??閿熻棄煤閿曞倸鐭楅柛鎰╁妿閺嗭箓鏌燂�??锟芥ɑ鍎曢柣鏃傚帶�???鍌炴煟閹炬娊顎楃紒銊ｅ劦濮婄粯鎷呴搹鐧告�??閿熶粙鏌涢幘瀵哥畾鐟滄壆濮电换娑虫嫹?閿熻姤顭囬惌瀣磼椤旇姤宕岋�??锟筋喖顭烽幃銏ゆ偂鎼达綆鍚嬮梻浣瑰劤濞存岸宕戦崨瀛樺仧闁哄啫鐗婇埛鎴︽偣閸ヮ亜鐨虹紒鐘冲哺閺岋繝宕ㄩ姘ｆ�?�閻庢鍠栭…鐑藉极閹剧粯鍋愰柟缁樺笩閳ь剙鐏濋�?�鍐Χ閸℃ê鏆楁繝娈垮枤閺屽宕愰幘顔解拻闁稿本鐟ㄩ崗�?勬煙閾忣偅宕岋拷?锟芥洜鏁诲浠嬵敇閻愭�??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖宕滆鐢盯鏌涳拷?锟筋煉锟???閿熶粙寮婚敓鐘茬闁靛ě鍐炬毇缂傚倷鐒﹂崝鏍�??锟芥繝鍥ц摕闁炽儲鍓氶崥�?�箹缁厜鍋撳畷鍥跺敹闂傚倷绶氶埀顒傚仜閼活垱鏅堕崜褏纾奸柣妯挎珪瀹曞矉锟???閿熺瓔鍠栭�?�閿嬩繆濮濆矈妲烽梺绋款儐閹瑰洭寮幇鏉跨＜婵炴垶鐟цぐ鍥╃磽閸屾瑨鍏屽┑�???娼ч悾婵堢矙濞嗙偓缍庢俊銈忕畳閿熴儲绂嶈ぐ鎺撶厵闁绘垶蓱閹牏绱掓潏鈺傛毄缂佽鲸鎸婚幏鍛村箵閹哄秴顥氭繝鐢靛仦閹稿宕洪崘顔肩；闁瑰墽绮敓锟???????闂備礁鐤囧Λ鍕�?囬悽鍛婃櫢闁跨噦�????闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???宕奸妷锔规嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵閸嬪嫭绂嶉敓锟???椤啴濡堕崱娆忣潷缂備緡鍠栧ù閿嬬珶閺囩喓闄勯柛娑橈功閸橆亝绻濋悽闈涗粶闁诲繑绻堝畷婵嬪箻椤旂晫鍘介梺瑙勫劤閸熷潡骞冮幋锔界厵濞撴艾鐏濇俊鐣岀磼缂佹绠烇�??锟芥洜鍠栭�?�锟??鎮欏▓鍨还闂傚倸鍊烽懗鍫曞箠閹捐搴婇柡灞诲劚缁犵�?鏌ㄩ悤鍌涘?濡ょ姷鍋涢崯鎾箖濠婂牊瀵犲璺虹焸閻涙捇姊绘担绋款棌闁绘挸鐗撳畷顖炲煛閸涱厾顓洪梺缁橆焽閺佹悂鏁嶅┑�?�拺缂佸瀵у﹢浼存煟閻�?潙濮傦拷?锟芥洘顨婇弫鎾绘晸閿燂拷??缂備浇椴哥敮锟狅�??锟藉璺哄窛妞ゆ挾濮冲鎾绘⒒閿燂拷?濞佳兾涘Δ鍛柈妞ゆ牗绮嶅畷鍙夌節闂堟侗鍎忛柣鎰躬閺屾洘寰勯崼婵堜患婵炲瓨绮嶉崕鎶芥箒闂佹寧绻傞幊搴ㄋ夎箛鏃傜閻忓繑鐗�?▍濠囨煙椤旇偐绉猴拷?锟芥洦鍋婂畷鐔碱敆娴ｇǹ澹嶉梻鍌欑閹芥粓宕戦幋锟??�?夐敓�????閸曘劉鍋撻弮鍫濈妞ゆ柨妲堣楠炴牗娼忛悙锟??�????闂佽法鍠曞Λ鍕綖閸ヮ剚鈷掑�?�姘ｅ亾婵炰匠鍥ㄥ亱闁糕剝銇傚☉銏╂晣闁绘柧�?�?ù鍕⒑閸愬弶鎯堥柟鍐茬箻閸╂盯骞嬮敂鐣屽幈闂婎偄娲﹂幐鎼佸箖閹达附鐓忛柛銉ｅ妿缁犳捇妫佹径�?�瘈濠电姴鍊归ˉ鐐电棯椤撱垻鐣洪柡宀嬬秮閺佹劙宕惰楠炲螖閻橀潧浠滄繛宸弮閵嗕礁顫滈�?顒勫箖閳哄拋鏁冮柨婵嗘矗缁ㄧ晫绱撻崒姘炬�??閿熶粙宕愭搴㈩偨闁跨喓濮寸壕濠氭煙閻戞﹩娈旈敓�????閸儲鐓熼柡鍌涱儥濞堢姵绻涢崗鑲╁ⅹ闁宠鍨块幃鈺嬫�??閿熺晫濮撮ˉ婵堢磼閻愵剙鍔ら柛姘儔楠炲牓濡搁妷顔藉缓闂佺硶鍓濋�?�鍛寸嵁鐎ｎ喗鈷戠紒瀣儥閸庢劙鏌熼悷鐗堝枠闁绘侗鍣ｅ浠嬪Ω閿燂�??椤庢捇姊洪崨濠勭細闁稿氦宕靛Σ鎰邦敋閳ь剙顫忕紒妯诲闁告縿鍎虫闂佽法鍣﹂敓锟???????濠电偠鎻徊浠嬪箹椤愇诲顫濋懜鐢靛幈闂佹寧妫侀褔鐛幇鐗堢厱閻庯綆鍋呭畷�?勬煙椤旀儳鍘达拷?锟筋喛娉涢埢搴ㄥ矗閵壯勶紡闂傚�?�鍊风欢姘焽閼姐�?�绶ら柛褎顧傛径鎰�?闁哄顕抽敃鍌涚厵闁绘鐗婄欢鑼磼閻樺啿鈻曢柡�???鍠撻�?顒傛暩鏋拷?锟芥繈姊洪柅鐐茶嫰婢т即鏌涳拷?锟筋煉锟???閿熶粙鐛�?崘銊ф殝闁归潧鍟块悧姘舵⒑閸涘﹤濮夐柛瀣崌閸┿垽宕奸妷锔兼嫹?閿熻姤绻涢崼婵堜虎闁哄鍠栭弻鐔碱敊閻撳簶鍋撻幖渚囨晪闁挎繂妫涢々鐑芥�?�閿濆懐浠涢柡鍜冪秮濮婅櫣绱掑Ο鑽ゅ弳闂佸湱鈷堥崑濠囨偘閿燂拷?楠炲洭鎮ч崼姘濠电偠鎻敓�????妞ゎ偄顦靛畷鎴︽偐缂佹鍘遍柟鍏兼儗閸犳牠鎮�?敂閿亾鐟欏嫭绀冩繛鑼枛�?�宕卞Δ濠傛�??????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閿燂�???闂佹寧绻傛鍛婃櫠娴煎瓨鐓熼柨鏇�?亾闁绘鎹囬獮鍐ㄎ旈崘鈺佹�?�闂佸憡娲﹂崜娑⑺囬妷鈺傗拺缂備焦顭囨晶顏堟煕濮橆剦鍎愮紒宀冮哺缁绘繈宕堕妸銉㈠亾婵犳碍鐓㈡俊顖滃皑缁辨岸鏌曟繛褍�?�弸鎴︽煥閻曞倹锟???闂佸憡娲﹂崑鍡涙偩濞差亝鈷戦柟绋挎捣缁犳挻绻涚仦鍌氬濠㈣娲樼粋鎺炴嫹?閿熺瓔鍋嗛崢閬嶆煟韫囨洖浠滃褌绮欓獮濠囧幢濡晲绨婚梺鍝勶�??锟介娆徫熼�?顒勬煥閻曞�?�锟???????婵＄偑鍊栭崝褏寰婇悾灞筋棜闁规儼濮ら埛鎴︽煕濠靛棗顏敓�????娴煎瓨鐓熼柍鍝勶工閻忥箓鏌曢崱鏇犵獢鐎殿喗鎸抽敓�????闁斥晛鍟悵鎶芥⒒娴ｈ鍋犻柛搴㈢矌娴狅箓骞嗚閻忓酣姊婚崒姘炬�??閿熶粙宕愰悜鑺ユ櫢闁跨噦�???????闂傚倷鑳舵灙妞ゆ垵妫濋獮鎰板箹娴ｅ湱鐣抽梻鍌欒兌缁垶鏁嬪┑鈽嗗灠閿曨亜鐣烽弴銏犵疀闁绘鐗忛崢浠嬫⒑鐟欏嫬鍔ら柣掳鍔庣划鍫嫹?閿熺瓔鍠楅悡娆愩亜閿燂拷?閺嬪鎳撻崸妤佺厵妞ゆ梻鏅幊鍥殽閻愬瓨宕屾鐐村浮�?�曞崬螣閾忚楔濠电姷鏁告慨鐢割敊閺嶎厼绐楁俊銈呭缂嶆﹢姊绘担鍛婂暈闁哄被鍔戦弻濠囨晲婢跺苯绁︽繝銏ｅ煐閸�?洜绮婚悷鎳婂綊鏁愰崶銊ユ畬婵炲瓨绮撴禍璺侯潖濞差亜绀堥柟缁樺笂缁ㄨ偐绱撴担绛嬪殭閻庢矮鍗抽獮鍐倻閽樺鎽曢梺闈涱檧閼靛綊骞忛搹鍦＝濞达絽澹婇崕蹇涙煟韫囨梻绠炴い銏☆殜閿燂拷?閹鸿櫕绂嶅⿰鍫熺厪濠电偛鐏濋崝婊勩亜閵壯冧户缂佽鲸甯掗悾婵嬪礃椤斿吋鎳欑紓鍌欒兌缁垳鎹㈤崼婵堟殾闁割偅娲嶉�?顒佺墵椤㈡牠顢楅�?�???煤閿曞�?�鍋傞柡鍥╁枔缁犻箖鏌燂�??锟芥绠撻柤绋跨秺閺屸槄�????閿熺瓔鍋嗛埊鏇犵磼缂佹娲达�??锟芥洩锟??????濠电姵顔栭崰鏍晝閵娿儮鏋嶉柨婵嗘处椤洟鏌熼悜妯烘闁绘梻鍎わ�??锟芥岸鏌＄仦璇插姷闁瑰嚖�????闂佽法鍠曟慨銈囨崲濠靛鍋ㄩ梻鍫熺◥閸濇鏌ｈ箛鎾剁闁荤啿鏅涢悾閿嬪閺夋垵鍞ㄩ悷婊勭矒�?�曠敻寮撮悙鈺傛杸闂佺粯锚绾绢參銆傞弻銉︾厱閻庯綆浜濋ˉ銏ゆ煛鐏炲墽銆掑ù鐙呯畵瀹曟粏顦俊鎻掔墦閺佹捇鏁撻敓锟????????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犲灚鍔栧瓭闂備緤�????閿熻棄鑻晶鍓х磼閻樿櫕灏柣锝囧厴�?�曞ジ寮撮妸锔芥珜闂備緤�????閿熻棄鑻晶鎵磼椤旂⒈鐓奸柟顔规櫇缁辨帒螣閻撳骸绠為梻鍌欑窔閳ь剚绋戝畵鍡樼箾娴ｅ啿娲ら崙鐘绘煟閺傚灝鎮戦柣鎾跺枛閺�?喖骞嗚閺嗛亶鏌￠崱娆忔灈闁哄瞼鍠栭幊鐘活敆婵犲啫锟????闂傚倷绀佹竟濠囧磻閸涱垱宕查柛鏇ㄥ�?�閸ヮ剦鏁囬柣鎰ㄦ櫆閿燂�??闂佽法鍣﹂敓�???????缂傚倸鍊搁崐鎼佹偋閸涘瓨鏅搁柨鐕傛嫹???濠碉紕鍋戦崐鏍ь啅婵犳艾纾婚柟鍓х帛閻撴洟鏌ｉ弬鎸庡暈缂傚秵鍨块弻锝夋晲婢跺鏆犵紓浣芥閺咁偆鍒掑▎蹇婃�?�闁绘劦鍓涚粔閬嶆⒒閸屾瑨鍏�?紒顕呭灡閻忔瑩鏌ｈ箛鎾剁闁荤噦濡囩划�?�吋閸℃鍤ら柣搴㈢⊕鑿ら柟椋庣帛缁绘稒娼忛崜褍鍩岄梺纭咁嚋缁绘繈鐛崱娑�?唶闁靛濡囬崢閬嶆⒑缂佹ɑ纾婚敓锟???娴ｅ湱顩插ù鐓庣摠閻撴瑦銇勯弬璇插婵炲眰鍊濋悰锟??�???閿涘嫮顔曢梺鐟邦嚟閸嬬喖骞婇崨�?�樼厱婵☆垵顕ч悘瀛樻叏婵犲啯銇濇鐐寸墵閹瑩骞撻幒鎳躲倝姊绘担鍛婂暈闁规瓕顕ч悾婵嬪箹娴ｅ摜鐣洪梺鐐藉劜閺嬬厧危閸儲鐓忛煫鍥ュ劤绾惧潡鏌涢敓锟???娴滆泛顫忓ú顏咁棃婵炴垼椴歌�?�闂備焦鎮堕崝宀勫箹椤愶箑鐓濓拷?锟姐儱顦婵嬫倵濞戞瑯鐒介柛妯绘�?�閺岋絾鎯旈婊呅ｉ梺绋款儏閹虫ǹ妫㈤梺鍓插亖閸庢煡鎮″☉銏★�??锟介柣鎰絻閳锋棃鏌嶉挊澶樻█闁硅棄鐖奸弫鎰緞鐎ｎ剙寮伴梻濠庡亜濞诧妇绮欓崼銉ョ；闁圭偓鏋煎Σ鍫熸叏濡櫣浜敓�????閸濆嫧鏀介柣妯虹仛閺嗏晠鏌涙惔銏犵仼鐎垫澘锕幐濠冪珶濠靛洦銇濆┑陇鍩栧鍕舵嫹?閿熺瓔鍋呴悵鏍ㄤ繆閻愵亷�????閿熺晫鎹㈤幇鐗堝亱闁糕剝鐟ф稉宥夋煛�?�ュ啫濡跨紒鐘荤畺閺屾盯鍩勯崘鐐暦缂備礁鍊搁澶愬蓟濞戙垺鍋勯梺鍨儏濞呫倝姊洪棃娑欐悙閻庢碍婢橀锝夘敋閳ь剙鐣烽幒鎴僵妞ゆ垼娉曠敮娑欑�?閻㈤潧袨闁搞劌顭烽獮濠囧箻缂佹ê浜遍梺绯曞墲缁嬫垿鎮￠敓锟???閺岀噦锟???閿熺晫枪娴犳粎绱掗悩闈涒枅婵﹨娅ｇ划娆撳礌閳╁啯鏆版俊鐐�??锟介崝灞轿涘┑�?�祦闁割偁鍎辨儫闂佸啿鎼崐鍛婄閾忓湱纾藉ù锝呭閸庢挻绻涙径瀣闁诡喗鍎崇叅妞ゅ繐鎳夐幏铏圭磽娴ｅ壊鍎愰悗绗涘喛鑰块柣�???鐗婇崣蹇斾繆椤栨簱瑙勬叏閸屾壕鍋撳▓鍨灍濠电偛锕顐�?礃椤旇偐锛滃┑鐐村灦閼瑰墽鏁ィ鍐┾拻濠电姴楠告禍婊勭箾鐏炲偊锟???閿熶粙銆�?弽顓炲窛闁哄鍨归崝�???顪冮妶鍡楃瑐闁绘帪濡囩划鍫ュ醇閵忋垻锛滃銈嗘煥閻忔繈宕ラ崷顓犵＜閺夊牄鍔岀粭鎺楁懚閿濆鏅搁柨鐕傛�??闂佸綊鍋婇崰姘枖閸ф鈷掗柛灞剧懅椤︼箓鏌熺喊鍗炰喊鐎规洦鍨堕�?�鏇㈡晝閳ь剛澹曡ぐ鎺撶厽闁绘梻枪椤ユ劙鏌★拷?锟筋亞效闁哄矉绻濆畷鍫曞Ψ閵壯傜棯闂備胶绮幐璇裁哄Ο鑽も攳濠电姴娴傞弫宥嗙�?婵犲倸鏆欏┑鈩冩そ濮婃椽宕妷銉︾亖闂佺ǹ顑囬崰鎾澄ｉ幇鏉跨闁哄啫鍊婚敍婊堟煥閻曞�?�锟?????婵犵數濮烽弫鎼佸磻閻旂厧鍌ㄧ憸蹇涘箲閵忕姈鐔兼惞鐟欏嫭顔曟繝鐢靛Т閿曘倕螞椤撶倣锝嗐偅閸愨晛浠╁┑顔矫晶鐣岀矙鐠囩潿搴ㄥ炊瑜濋煬顒勬煙椤旂晫鎳囨い銏℃瀹曠喖濡搁妷銈咁棜闂備線娼ч悧鍡浰囬婊冾棜濠电姵纰嶉悡鏇㈡煛閸ャ儱濡奸柣搴墴閺屾盯濡烽敐鍛�?�缂傚�?�绉村ú顓㈠蓟閺囩喓绠剧憸宥夊嫉椤掑嫭鐓ラ柕鍫濐槹閳锋帒霉閿濆懏鎲哥紒澶屽劋娣囧﹪顢曢�?鈥充淮闂佽鍠氶崑銈夊极閸愵喖纾兼慨妯诲敾缁遍亶姊婚敓锟???濞佳嗗闂佸搫鎳忕划鎾诲箖閿熺姴鍗抽柣鏃囨椤旀洟姊洪悷閭﹀殶闁稿孩鍨垮畷妤咁敆閸曨剛鍘遍梺鍝勫暙閸婃悂寮稿☉銏＄厸閻忕偛澧介埥澶愭懚閿濆鐓曢煫鍥ㄦ尭閹垶鎱ㄩ敐鍛闁宠鍨块、娆戞兜闁垮鏆版繝纰夌磿閸嬬姴螞閸曨垱鍋╅柣鎴ｆ鎯熼梺鎸庢煥婢т粙鎯侀崼銉︹拺闁告稑锕ユ径鍕煕閹惧鎳冮柍璇茬Ч楠炲鎮欓幍顔剧暰闂佽法鍣﹂敓�?????????闂傚倸鍊搁崐闈╂�??閿熺瓔鍓涢埀顒佸嚬閸樺墽鍒掗埡鍛亜闁绘挸楠搁懓鍨攽閳藉棗鐏ｉ柍宄扮墕鐓ら柟闂寸劍閳锋垹鎲搁悧鍫濈瑲闁挎稓鍠栭弻锝夊箳閻愮數鏆ら悗娈垮枟瑜板啴銈导鏉戝窛妞ゆ牗绮ｇ槐鍙夌�?閻㈤潧浠﹂柛銊ョ埣閺佸啴鍩￠崨顓狅紵闂佸綊鍋婇崢瑙勭濠婂牊鏅搁柨鐕傛嫹??婵犵妲呴崑鍕疮椤愶讣缍栭煫鍥ㄧ⊕閹偤鏌涢敂璇插箻闁挎稒绮岄埞鎴�?煡閸℃浠╅梺鍦拡閸嬪﹪鏁愰悙宸悑闁告侗浜濋敓锟???闂備胶绮崝鏍亹閸愵喖绠栭柟杈鹃檮閻撶喖鏌ｉ敓�????缁诲倿骞婃惔銊ュ瀭婵犻潧娲㈡禍婊堟煙閹冭埞闁诲繆鏅濈槐鎺楁偐閻戞褰ф繛锝呮搐閿曨亝淇婇崼鏇炵妞ゆ挾鍋涢�?�澶愭⒒娴ｈ鍋犻柛濠冩礋钘濋梻鍫熶緱濞兼牗绻涘顔荤盎濞磋偐锟??閺屾盯寮撮妸銉ョ闂佸搫顑呭Λ婵嗩潖閾忚瀚氶柤纰卞墰椤斿姊洪崨濠冣拹闁挎洏鍨烘穱濠囨偨缁嬭法锟??闂佸搫顦冲▔鏇㈩敊婵犲洦鈷戦悷娆忓閸斻倝鏌ｆ幊閸旀垿骞冮悽绋跨婵炴潙顑嗛敓锟???闂備胶绮敃鈺呭窗閺嶎厽鍊堕弶鍫涘妿缁犳儳顭跨捄渚剳婵炴彃鐡ㄩ妵鍕閿涘嫬鈷岄悗瑙勬�?瀹曨剟鍩ユ径濞㈢喖寮拌箛鏇炲絺闂傚�?�鍊烽懗鍓佸垝椤栫儑�????閿熶粙宕堕埡浣哥亰濡炪�?�鐗滈崑娑㈡偂閺囥垺鐓欓弶鍫ョ畺濡绢噣鏌ｉ幘瀛樼缂佺粯绻堝Λ鍐ㄢ槈濮�?棔鎮ｉ梻浣告啞濮婂綊鎳濇ィ鍐╃畳闂備胶绮敋缁剧虎鍙冮幆�?嬫嫹?閿熺瓔鍠楅悡蹇涙煕閵夋垵鍠氭导鍐⒑鏉炴壆顦﹂柛鐔告綑閻ｇ兘骞掗幋锟??顫嶅┑鐐叉閹稿寮冲Ο琛℃斀闁挎稑�?�禍濂告煕婵炲尅锟???閿熻棄鐣烽幋�???�?嬫い鎾跺枎鎼村﹪姊洪崷顓炲妺婵﹤缍婇敐鐐哄即閵忥紕鍘甸梺缁樺灦閿氭繛鍫ョ畺閺岋綁寮�?崒姘�?闁诲孩纰嶉悢顒勫箯閿燂�???闂佽法鍠曞Λ鍕珶婵犲洤绐楅柟鐑橆殔绾惧鏌熼幑鎰靛殭缂佺姾宕电槐鎾存媴妤犮劍�?搁獮蹇撁洪鍛嫼闂佸憡绋戦敃锕傚煡婢舵劖鐓ラ柡鍥朵簻椤╊剛绱掓潏銊�?碍妞ゎ偅绻堥幊婊堟偨闂堟稑绠為梻浣烘�?閸氬鎮鹃鍫濈９闁哄稁鍘介崑鐔搞亜韫囨挻鍣峰ù婊勭矒閺屾洘绻濊箛鎿冩喘闂佺懓鍟块崯鎾蓟瀹ュ洦鍠嗛柛鏇ㄥ亞娴煎矂姊烘潪鎵槮缂佸鎳撻悾鐑芥偄绾拌鲸鏅濋梺鏂ユ櫅閸燁垳娆㈠鑸碘拻闁稿本鐟ㄩ崗宀勫几椤忓牊鐓ラ柡鍥崝锔兼�??閿熻姤娲栫紞濠傜暦瑜版帩鏁婇柣鎰靛墯椤旀洟姊绘担鍛婃儓婵炲眰鍨藉畷纭呫亹閹烘挸鐝旈梺缁樻煥閸氬鎮¤箛鎿冪唵閻犻缚娅ｆ晶鏇㈡煕閺備紮锟???閿熶粙濡甸崟顖氭婵炲棛鍋撻埢鍫濃攽椤旂》鏀绘俊鐐扮矙閻涱噣寮介鐕傛嫹?閿熶粙鏌熺紒妯虹瑨閾绘岸姊婚崒娆戭槮闁规祴鍓濈粭鐔肺旈崨顓犵崶濠德帮�??锟介幏�?�极婵犲洦鐓涢柛銉㈡櫅閺嬫棃鏌ㄩ悤鍌涘�??闂佽楠搁敓�????闁告濞婂銊╁�?閻戝棛鍞甸梺璺ㄥ櫐閿燂拷??闂佽法鍣﹂敓�?????婵＄偑鍊栫敮濠勭矆娴ｈ鍙忥�??锟姐儱绻戦敓�?????闂佽法鍠曟慨銈吤洪敓�????瀹曞綊宕稿Δ鍐ㄧウ濠碘槅鍨伴幊娆愭償椤垶鏅為柣鐘充航閸斿骸鈻旈崹顔规�?闁挎稑�?�禍濂告煕婵犲啰澧碉拷?锟芥洘绻嗛ˇ杈炬嫹?閿熻姤婢�?敃顏勭暦缁嬭锟??鎷呯粙鍨棗闂傚倷绀佸﹢閬嶅磿閵堝�????閿熶粙宕卞☉娆忎簵闂�?潧顦弲婊堟偂閻斿吋鏅搁柨鐕傛嫹??????????濠电姷鏁告慨鐑斤�??锟介鐐潟闁哄洢鍨圭壕濠氭煙鏉堝墽鐣辩痪鎯х秺閺岋拷?锟界暤椤旇壈瀚伴柡鍛У缁绘繈鎮介棃娴讹綁鏌ら悷鏉库挃濠㈣娲樼换婵嗩潩椤撶姴骞嶉梻浣虹帛閸旓箓宕滃☉銏犳辈婵☆垰銈介悷鎵冲牚闁告洦鍘鹃悡澶愭⒑閸濆嫮鐒跨紒缁樼箓閻ｇ兘宕奸弴鐐茬彉闂佹眹鍨归悘姘跺疾閼测晝纾介柛灞剧懅椤︼附銇勯敂璺ㄧ煓鐎规洘婢樿灃闁告侗鍘欓敃鍌涚厱闁哄洢鍔岄悘鐘炽亜椤愩垺鍤囬柡灞界Ч閸┾剝鎷呴崨濠冾�?婵＄偑鍊х紓姘跺础閸愬樊娼栭柣鎴炆戞慨婊堟煙濞堝灝娅樻俊宸櫍濮婃椽宕妷銉︼�??锟介梺鍦�?归崯鍧楁偩�?�勬噴娲敂閸曨厼濮︽俊鐐�??锟界敮濠囨⒔瀹ュ棛顩叉繝濠傜墛閻撴瑩鏌ｉ幋鐏活亪鎮橀妷鈺傜厓鐟滄粓宕滃☉姘灊妞ゆ牗绮庨惌娆忣熆鐠鸿�?鐪嬮柛姘儏椤法鎹勬笟顖氬壋闂佸憡顭囬崑鎾舵崲濠靛棌鏋旈柛顭戝枟閻忓秹姊洪崨濠冣拹婵炶尙鍠栭弫鎾绘晸閿燂拷??婵＄偑鍊栫敮濠勬閳ユ枼鏋旀俊顖欒閻斿棝鎮峰▎蹇擃仾閿燂拷?鐎ｎ喗鐓欑紒瀣皡锟??鑽ょ磼閺冨�?�鏋庨柍瑙勫灴�?�曞崬鈻庨幊韬插姂濮婄儤娼幍顔煎闂佸憡姊归悷銉╂偩閻戠瓔鏁傞柛娑卞枛椤庢捇姊洪棃鈺佺槣闁告﹢绠栭崺銉�?緞婵炵偓�???闂佹寧绋戯拷?锟筋剚绂嶆總鍛婄厱濠电姴鍟粈鍫ユ煙楠炲灝鐏叉鐐叉喘椤㈡瑩鎮锋０浣割棜??闂備焦鎮堕崕婊堝礃閵婏富鍚囬梻鍌氾拷?锟界粈锟??骞栭锟??鐤柣妯款嚙绾惧鏌熼幆褏鍘旈幖娣妼閻愬﹦鎲稿┑�?�彆妞ゆ巻鍋撻柍瑙勫灴閸ㄦ儳鐣烽崶褏鍘介柣搴ゎ潐濞叉鏁幒妤嬬稏婵犻潧顑愰弫鍐煏韫囧﹥娅嗘い銉節濮婂宕掑顑藉亾閹间礁纾瑰�?�捣閻棝鏌ㄩ悤鍌涘?闂佽鍠栧鈥崇暦閸洦鏁嗗┑鐘插閳笺倕鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪即閵忕姴鐎梺绋跨灱閸嬬偤鎮￠弴鐘冲枑閹兼番鍔屾濠电姴锕ら悧鍡涙倿閸偁浜滈柟杈剧稻绾埖銇勯敂鑲╃暤闁哄苯绉堕幏鐘诲蓟閵夈儱鍙婃俊銈囧Х閸嬬偤鏁冮姀銈呯鐟滅増甯╅弫鍐┿亜閹板墎绉垫俊顐犲姂濮婂宕掑顑藉亾妞嬪孩顐芥慨姗嗗墻閻掔晫鎲搁弮鍫濈畺鐟滄柨鐣烽崡鐐╂瀻閻忕偞鍨濇竟鏇炩攽椤旂瓔鐒介柛妯犲洤鍑犻柣鏂挎憸缁犻箖鏌ｉ幘鍐茬槰闁绘捁鍋愰埀顒侇問閸ｎ噣宕抽敐鍛殾濠靛倸鎲￠崑鍕煕濞嗗浚妲告い蹇曞劋缁绘繈鎮介棃娑楀摋闂佽妞挎禍鐐差嚗婵犲啰顩烽悗锝庝簽閻ゅ懘姊虹捄銊ユ灁濠殿喗鎸抽幃鍧楊敋閳ь剟寮婚敐澶婄�?妞ゆ梻鍘ф俊娲⒑缂佹ɑ灏伴柣鐔濆懏顫曢柟铏瑰仦閿燂�???闂佽法鍠撻悺鏃堝磻閹烘纾块柕澶嗘櫆閻撶喖鏌熼崜褍浠洪柛瀣ㄥ灲閺岋拷?锟界暆閳ь剟宕伴弽顓ㄦ�??閿熻棄鈻庨幘宕囩暰閻熸粌绉归悰顕嗘嫹?閿熺瓔鍠楅埛鎴﹀级閻愭潙顥嬫い锔肩畵閺屾稒绻濋崒娑樹淮濡ょ姷鍋涢崯顐�?煝鎼淬劌绠奸柛鎰ㄦ櫆濞呭矂姊婚敓�????閳ь剛鍋涢懟顖涙櫠椤栫偞鐓欐い鏍ㄧ⊕閳锋劗绱掔紒妯肩疄鐎规洘甯掕灃濞达�?顫夊鎴︽⒒閸屾瑨鍏�?紒顕呭灦瀹曟繈寮借閻掕姤绻涢崱妯诲鞍闁稿﹤鐖奸弻锝夊棘閸喗鍊梺缁樻尰濞茬喖寮婚弴鐔虹闁割煈鍠栨慨銏㈢磽娴ｅ壊妲规俊鐐扮矙瀵鎮㈢喊杈ㄦ櫓闂佷紮绲介張顒勫闯椤撶姷纾藉ù锝堟鐢稓绱掔拠鑼闁伙絿鍏橀弫鎾绘晸閿燂�???闂佽桨绀�?崐濠氬箲閸曨垰惟鐟滃酣寮查妸鈺傗拻闁稿本鑹鹃�?顒傚厴閹虫宕奸弴鐐电枃闂佽宕�?褏绮荤憴鍕�?簻闁规壋鏅涢�?顒侇殜閹矂骞樼紒妯煎幗闂佺鎻徊楣兯夋径鎰櫢闁跨噦�????????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕節閻㈤潧校妞ゆ梹鐗犲畷鏉课旈崨顓囷附绻涢幋娆忕仼缁炬儳顭烽弻鐔煎箲閹邦啩婊堟煟閻旂ǹ顥愰柛顐邯閺屾盯鍩勯崘鍓у姺闂侀潧妫欓崝鏇�??锟介崘顔嘉ч幖杈炬�??閿熺晫鐩庣紓鍌欒兌缁垶宕濆Δ鍛煑闁告侗鍙庡〒濠氭煏閸繃鍣界紒鐘卞嵆閹顫濋梻�?�告晼濠碉拷?锟藉级閸�?瑥鐣锋總绋垮嵆闁绘柨寮讹�??锟藉ジ姊绘担鍛婂暈缂佸鍨块弫鍐Ψ閿燂拷?缁剁偤鏌涢弴銊ョ仭闁绘挻娲樻穱濠囶敍濠靛棗鎯為梺娲诲幗鐢繝寮婚悢纰辨晩閻熸瑥�?�悵鏍磽娴ｄ粙鍝洪悽顖涘笩閻忔帡姊虹紒妯诲碍濡ょ姴鎽滅划濠氭倷鐎靛摜鐦堥梺姹囧灲濞佳冩毄闂備浇妗ㄧ粈�???骞夐敓鐘茬疄闁靛ň鏅涚粻缁樸亜閺冨洤浜归柡灞界墕椤啴濡堕崱娆忣潷缂備緡鍠栭柊锝夊箚锟??鍕耿婵炴垶鐟ч崢閬嶆⒑闁稑宓嗘繛浣冲洤鍑犻柣鏂垮悑閻撶喖鏌熼幆褜鍤熸繛鍙夋尦閺岋紕浠﹂崜褉妲堥梺�?�犳椤﹂潧鐣烽敓鐘筹拷?锟介柤纰卞墻閸熷姊婚崒娆掑厡缁绢厼鐖煎鏌ヮ敂閸℃绛忛梺绉嗗嫷娈旈柣鎺戠仛閵囧嫰骞掑鍥獥闂佸摜鍠庣换�???寮诲☉銏″亹鐎规洖娲ら敓�???????闂傚倸鍊风粈�???鎮樺┑�?�垫晞闁告洦鍘藉畷鏌ユ煕閳╁啰鈯曢柣鎾跺枛閺�?喐娼忛崜褍鍩岄悶姘哺濮婃椽宕崟锟??娅ら梺璇″枛閸婂灝顕ｆ繝姘╅柍鍝勶�??锟芥禍鐐烘煥閻曞倹锟???????闂傚倸鍊搁崐鎼佸磹妞嬪孩顐芥慨妯挎硾閻掑灚銇勯幒鎴�??閿熻姤绂掑⿰鍫熺厾婵炶尪顕ч悘锟犳煥閻曞�?�锟?????闂備礁鎼惌澶岀礊閳ь剛绱掗悩宕囨创鐎殿噮鍓熷畷褰掝敊閼恒儱娈樻繝寰峰府锟???閿熻姤鎱ㄩ悜钘夌；婵炴垯鍨洪崑�?�煙閸撗呯瘈缂佽妫濋弻鐔兼⒒鐎靛壊妲�?柛鐑嗗灠椤啴濡堕崱姗嗘⒖濠碘槅鍋勶�??锟筋喚妲愰幘璇茬缂備焦菤閹风粯绻涙潏鍓хК婵炲拑缍佹俊瀛樼�?閸ャ劎鍘遍梺瑙勫劤椤曨厾绮婚悙鐑樼厪闁糕剝顨呴弳锝忔�??閿熻姤娲忛崝宥咁焽韫囨稑�?堢憸蹇涘煟閵堝棔绻嗛柣鎰典簻閳ь剚鐗犲畷婵嬪箣閿燂�??绾捐淇婇妶鍛殭妞ゃ儲�?搁弻�???螣娓氼垱锛嗛悷婊呭鐢寮查弻銉︾厱婵炴垵宕鐐繆椤愩垼�?�伴柍瑙勫灴濡鹃亶鎮樿箛锝勯偗闁挎繄鍋炲鍕舵嫹?閿熺瓔鍏�?弨铏節閻㈤潧孝婵炶绠撳畷鎰版倻閼恒儳鍘靛┑鐐茬墕閻忔繈寮搁妶澶嬬厽闁规儳鐡ㄥ畷宀勬煙椤旂瓔娈旈柍缁樻崌�?�曞綊顢欓悾灞奸偗濠碉紕鍋戦崐銈夊储妤ｅ啫绀傛俊顖欒閸ゆ洘銇勯幇鈺佺労闁告艾顑呴�?�璺ㄦ崉閻氭潙濮涘銈忛檮濠㈡﹢鈥旈崘顔嘉ч柛娑卞灣椤斿洭姊洪悷鏉挎毐閻庢稈鏅犲畷姘�?閸愵煈鍤ら柣搴㈢⊕鑿ら柟閿嬫そ濮婃椽鎮℃惔顔界稐闂佺ǹ锕ュú鏍偤椤撶喓�???闁汇垽娼ф禒鈺傘亜閺囩喓鐭�?紒顔碱煼楠炴帒螖閳ь剚顢婇梻浣告贡婢ф顭垮Ο鑲╃焼闁告劏鏂傛禍婊堟煛閸モ晛浠︽い銉уХ缁辨帪�????閿熺瓔浜炵粻缁樻叏婵犲啯銇濇鐐寸墵閹瑩骞撻幒鎳躲倝姊绘担鍛婂暈闁规瓕顕ч悾婵嬪箹娴ｅ憡妲┑鐐村灟閸ㄥ湱绮婚敐澶嬬叆闁哄啫娲﹂ˉ澶娒归敓�????閸ㄨ泛顫忓ú顏勭闁绘劖褰冩慨椋庣磽娴ｇǹ绾ф俊鐐舵閻ｇ兘骞嬮敓�????缁犺崵绱撴担鑲℃垿宕曢鍕垫富闁靛牆妫楁慨鍌炴煕婵犲啯灏甸柤娲憾楠炴﹢顢欑憴锝嗗闂備胶枪閺堫剟鎮疯瀹曟繂顓兼径瀣幍濡炪�?�妫�?崑鎰板春閿濆洠鍋撶憴鍕缂佽妫涚划璇测槈閵忕姷顔掗梺褰掑亰閸樻儳煤鐎电硶鍋撶憴鍕闁哥姵鐗犻妴浣糕槈濡攱顫嶅┑鈽嗗灥椤宕戦崨瀛樷拻闁稿本鐟ㄩ崗锟??绱掗鍛仸鐎规洖缍婇幃锟犵嵁椤掍胶娲达�??锟芥洜鍠栭弫鎾绘晸閿燂拷??闂佸憡姊瑰Λ鍐潖婵犳艾纾兼繛鍡樺灥婵′粙鏌ｆ惔锝囨嚄闁搞儜鍡樻啺闂備線娼чオ鐢告⒔閸曨�?鏋嶉柣妯款梿瑜版帗鍋愶拷?锟藉壊鍠栭崜閬嶆⒑缁嬪潡顎楅柨鏇ㄤ邯瀵鈽夐姀鈺傛櫇闂佺粯蓱瑜板啯鎱ㄩ弴銏�?拺闁规儼濮ら弫閬嶆煕閵娿儲鍋ワ拷?锟筋喛顕ч埥澶娢熼柨�?�垫綌婵犳鍠楅〃鍛存偋婵犲洤鏋�?柣鎰靛墰閿燂�??闂侀潧楠忕徊鍓ф兜妤ｅ啯鍊垫慨妯煎帶婢у瓨绻濋埀顒佹媴缁洘�???闂佺粯枪椤曟粌顔忛妷鈺傜厵闁告劖褰冮銏㈢磼閸屾稑绗╂い�???寮堕妵鍕敇閳╁啰銆婇梺鐟板级閹稿啿鐣烽悢纰辨晢闁稿被鍊栨晥闂備浇顕у锕傦綖婢舵劖鏅搁柨鐕傛�???闂備礁澧界划顖炴偋閺囥垺绠掗梻浣瑰缁诲倿骞婃惔锝囨／鐟滄棃骞冮敓锟???椤繈顢曢妶鍥╁幆婵犳鍠栭敃锔惧垝椤栫偛绠柛娑欐綑�?�告繈姊婚崼鐔猴�??锟界紒澶庢閳ь剚顔栭崰姘跺极婵犳熬锟???閿熻棄螖閸涱厾顦伴梺璺ㄥ櫐閿燂拷??婵炲濯崣鍐潖濞差亝顥堟繛娣�?劚閻楁挸顕ｉ幓鎺嗘婵ǹ浜悞濂告⒑缁嬫寧婀板瑙勬礋�?�曟垿骞樼拠鑼槯婵犮垼娉涢敃锝嗙珶閺囥垺鈷掑ù锝呮啞閸熺偞绻涚拠褏鐣碉拷?锟芥洘绮岄埥澶愬閻樻彃浜堕梻浣圭湽閸ㄥ綊骞夐敓鐘茬厱闁硅揪闄勯悡娆愩亜閺嵮勵棞閻庢凹鍣ｉ妴鍛鐎涙ǚ鎷虹紓浣割儐椤戞瑩宕曡箛娑欑厵闁告劖鐓￠崣鍕煙椤旇棄鍔ら柣锝忕節楠炲秹顢欓懞銉ф殾闂傚倷绶氶埀顒傚仜閼活垱鏅堕敓锟?????濠碉紕鍋戦崐鏍暜閹烘绐楁慨姗嗗墻閻掍粙鏌熼柇�???骞樼紒鐘荤畺閺屾稑鈻庤箛锝嗭�??锟介梺鍏兼緲濞硷繝寮婚悢纰辨晪闁糕剝鐟ч惁鍫ユ⒑閹肩偛濮傜紒鐘崇墵閻涱噣宕堕妸�???顎撻梺鍛婄☉楗挳宕ュ▎鎰瘈闁汇垽娼у暩闂佽桨绀�?幉锟犲箞閵娾晜鍋ㄩ柛娑橈工濞堢偤姊虹拠鈥筹拷?锟介柛鏇ㄥ墯椤斿洭姊婚崒姘炬�??閿熶粙宕愭搴㈩偨婵﹩鍓﹂悞鐣屾喐閺冨洦顥ゆ俊鐐�??锟介幐鍫曞垂閸︻厼顥氶柛褎顨嗛悡娆撴煙椤栨粌顣兼い銉ヮ槸闇夐柤娴嬫櫅閳诲牊顨ラ悙瀵稿ⅹ閼挎劙鏌ㄩ悤鍌涘?婵犵锟???閿熺晫鐭欓柡灞界Ч閺岊煉锟???閿熺瓔浜為悷銊╂⒒閸パ屾█闁哄被鍔岄埞鎴�?幢濡儤顏￠梻浣告憸閸犳捇宕戦妶澶婅摕闁绘梻鈷堥弫宥嗘叏濡搫鑸归柍顏嗘暬濮婅櫣鎷犻垾铏仌濠电偛顦伴惄顖炴晲閻愭祴�?介悗锝庡亜娴滄鏌熼悡搴ｆ憼缂佽鍊垮鎼佸醇閵夛妇鍘介柟鍏肩暘閸娿倕顭囬幇顓犵闁告瑥顥㈤鍡�?疾闂備胶绮濠氬储瑜旈幏鎴︽偄閸忚偐鍘遍梺鏂ユ櫅閸犳艾鈻撻�?銈嗙厱婵﹩鍓﹂崕鏃堟煛鐏炲墽鈽夐柍钘夘�?瀹曪繝鎮欓懠顒夊晪闂傚�?�绶氶埀顒傚仜閼活垱鏅舵繝姘厱婵炲棗绻愰弳娆愩亜椤愩垻绠婚柟鐓庣秺瀹曠兘顢�?悩闈涘箚闂傚倷绀佸﹢杈ㄧ仚闁诲孩绋堥弲鐘荤嵁韫囨梹缍囬柍鍝勫暟閿涙繃绻涢幘纾嬪婵炲眰鍊濆绋库槈濮樿京锛滄繝銏ｆ硾閺堫剟宕甸埀顒勬⒑娴兼瑧绉敓锟???鏉堚斁鍋撻棃娑栧仮鐎殿喖鐖奸獮�?�偐閸偅绶梻鍌氾拷?锟介懗鍓佸垝椤栫儑锟???閿熶粙宕拷?锟芥ê浜遍棅顐㈡处缁嬫垿宕掗妸銉冨綊鎮╁顔煎壉闂佹娊�?遍崹鍧楀箖瑜版帒绠掗柟鐑樺灥椤牆鈹戦悙鍙夊櫤闁告梹鐟╁濠氭偄閻撳海顦╅梺闈涚墕濡顢旈敓锟????闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛鎾茬閸ㄦ繃銇勯弽顐㈠壋闁瑰嚖�????闂佽法鍠嶇划娆忕暦閵娾晩鏁囬柛銉ｅ妿閳藉鏌嶉挊澶樻Ц妞ゎ偅绻堥弫鎾绘晸閿燂拷??闂佽绻愰敃銈夛�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡奸敓锟???鏉堚晛鍨濆┑鐘崇閹偞銇勯幇鍓佺？缂佺姵宀稿娲濞戞艾顣洪柣搴㈠嚬閸ㄨ泛鐣烽敓�????閻ｆ繈宕熼鍌氬�???濠电偛鐡ㄧ划�?勬偉閻撳寒鍤曞┑鐘崇閺呮煡鏌涢鐘茬伄闁哄鎮傚娲传閸曨剙绐涢梺绋款儐閿曘垹鐣烽锔芥櫢闁跨噦�????濡炪値浜滈崯瀛樹繆閸洖骞㈡俊顖氱仢娴滄牠姊绘担鍛婂暈婵炶闄勭粋宥夋�?�閻㈠吀绗夊┑顔斤供閸樺墽寮ч�?顒勬煥閻曞�?�锟???????闂傚倷鑳堕�?�濠囶敋濠婂懏宕叉繝闈涱儏缁犳牠鏌ㄩ悢鍝勑㈤敓锟???閸愨斂浜滈柡鍐ㄦ处椤ュ霉閿燂拷?閸樺ジ鍩為幋锔斤�??锟介柛娆忣樈濡偟绱撴担铏瑰笡闁告梹鐟╅妴锟??寮崼婵堝幐闂佸憡渚楅崰姘跺储娴犲鏅搁柨鐕傛嫹????闂佽绻愭蹇曠不閹剧粯鏅搁柨鐕傛嫹???闂備礁鎽滄慨鐢告偋閻樿违濞达絿纭堕弸搴ㄦ煙鐎电ǹ浠滈柡�?��??锟藉娲川婵犲啫顦╅梺鍛婃尰缁嬫牠濡甸幇鏉垮窛閻庢稒菤閹风粯绻涙潏鍓хМ妞ゃ儲鎸荤粙澶愭嚑椤掑倻锛滈梺鍦帛鐢宕戦妷褉鍋撶憴鍕妞ゃ劌鎳撻悘鎺楁⒑閹呯妞ゎ偄顦埢鎾淬偅閸愨斁鎷洪梺鍛婃尰瑜板啯绂嶅┑鍥╃闁告瑥锟??閼板尅锟???閿熻姤娲滈�?�锟??骞忛敓锟????闂佽法鍠撻悺鏃堝窗濡ゅ懏鍋傞柡鍥╁枂娴滄粍銇勯幘璺烘瀻闁诲繈鍎遍湁婵犲ň鍋撶紒顔界懇�?�鈽夐姀鈥充簻闂備礁鐏濋鍛村几閻樻祴鏀芥い鏃傦�??锟藉銉︺亜椤撶偛妲婚柣锝囧厴楠炴帡骞嬮鐔峰厞婵＄偑鍊栭崹鐓幬涢崟顒傤洸闁诡垎灞惧瘜闁诲函缍嗘禍婵嬪箲閿濆鐓熸い鎾跺仦椤ユ粓鏌曢崱妯虹瑨妞ゎ偅绻堥弫鎰板川閿燂拷?椤ユ艾鈹戞幊閸婃鎱ㄩ悜钘夌；闁绘劗鍎ら崑�?�煟濡湱涓查柟鍑ゆ嫹?闂佽法鍠嶇划娆忣嚕閹绢喖顫呴柍鈺佸暞閻濇牠姊婚敓�????閳ь剛鍋涢懟顖涙櫠閹殿喚纾兼い鏃傗拡閻撳ジ鏌熼瑙勬珚闁圭绻濇俊鍫曞川椤撶姴顕遍梻鍌氾拷?锟介悞锕傚箖閸洖纾挎い鏍仜锟??澶愬箹濞ｎ剙濡奸柣鎿勬嫹?閿熺瓔鐔嗛悹楦挎閻忚京鐥幆褋鍋㈤柡宀嬬到铻ｉ柧蹇曟缁辩偞绻濋敓�????閸涱喗姣堥梺鍝勭焿缁辨洘绂掗敃鍌氱鐟滃危閸儲鈷戝ù鍏肩懅缁嬪鏌ㄩ悤鍌涘�????濠碉紕鍋戦崐鏍暜閹烘柡鍋撳鐓庡濠㈣娲滅槐鎺懳熼懖鈺婂晭闂備胶鎳撻悺銊╂偡閵夆晜鍊舵い蹇撶墛閸婂灚鎱ㄥ鍡�?闁搞�?�娲弻鈥崇暆鐎ｎ剛袦閻庢鍣崜鐔风暦瑜版帩鏁婇柡鍌橈�??锟介敓锟????闂佽法鍠嶇划娆忣潖閾忓湱纾兼俊顖濐嚙閽勫ジ姊虹粙鎸庢崳闁轰浇顕ч锝嗙�?濮橆厽娅滄繝銏ｆ硾閿曘儵藟濠靛鈷戦柛锔诲帎閸︻厸鍋撳☉鎺撴珚鐎规洘娲熼獮妯肩磼濡�?鍋撻崹顐ょ闁瑰鍋熼幊鍛磼閻樻剚鐒界紒杈ㄥ笚濞煎繘濡搁妷锕佺檨闂備浇顕栭崰妤呮偡閳哄拑锟???閿熻棄螖閸涱厾鍔�?銈嗗笒鐎氼剛绮堟径鎰厪闁割偅绻嶅Σ褰掓煟閹惧瓨�?冮柟渚垮妼椤粓宕遍敓锟???閳锋帡姊虹粙鍨劉婵﹤缍婇妴鍐Ψ閳哄偊�????閿熶粙鏌ょ喊鍗炲闁愁亜鐏氱换婵堝枈濡搫鈷夐梺璇�?�枛閸婅绌辨繝鍥ㄧ叆閻庯綆鍋勯崝鍛存⒑闂堟稓绠氭俊鎻掓噹铻為柛鎰靛枟閳锋垹绱掗娑欑闁哄缍婇弻娑虫�??閿熺瓔鍋呯亸顓熴亜椤忓嫬鏆ｅ┑鈥崇埣瀹曞崬螖閸愵亝鍣梻浣筋嚙鐎涒晠宕欒ぐ鎺戠煑闁告劑鍔庨敓�????????婵＄偑鍊曠换瀣倿閿曞�?�鏅搁柨鐕傛�??闂傚倸鍊烽懗鍓佸垝椤栨繃鎳岄柣鐔哥矋濠㈡﹢宕幘顕嗘�??閿熶粙寮�?崼婢冾熆鐠轰警鍎戦柛姗堟嫹???婵＄偑鍊栭崝褏寰婇悾灞芥瀳鐎广儱鎷嬪〒濠氭煏閸繈顎�?ù婊勭箘缁辨帞鎷犻懠锟??鈪靛Δ鐘靛仜閸燁偊鍩㈡惔銊ョ闁告劏鏅滃▍�?勬⒒閿燂�??閳ь剛鍋涢懟顖涙櫠鐎涙ǜ浜滈柕蹇婂墲椤ュ牓鏌ㄩ悤鍌涘�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕闈涱潖婵犳艾纾兼繛鍡樺笒閿燂�???闂傚倷鐒︼拷?锟窖兠鸿箛娑樼９婵犻潧顑呴悘鎶芥煥閻曞�?�锟???闂佷紮缍囩换婵嬪蓟閸ヮ剚鏅搁柨鐕傛嫹?濠电偛鐗勯崝鎴濐潖閾忚鍠嗛柛鏇ㄥ亜婵憡绻濆▓鍨灁闁稿﹥绻傞锝夊箵閹哄棗鐗氶梺鍓插亞閸犳捇宕㈡禒�?�拺闁圭ǹ娴风粻鎾绘煙閾忣偄濮嶉柟顔斤�?�閺屽棗顓奸崱娆忓箺??闂備胶绮�?�鍛存晝閿曞倸绠查柕蹇曞Л�???浠嬫倵閿濆骸浜滃ù鐘虫そ濮婂宕掑鍗烆杸闂佽法鍣﹂敓�?????闂備線娼х换鍫ュ磹閺嶎厽鍋傞柡鍥╁亹锟??浠嬫煟濡绲婚柡鍡欏仱閺佹捇鏁撻敓�?????????婵＄偑鍊栧Λ浣规叏閵堝纾归柟閭﹀厴锟??浠嬫⒔閸ヮ剙鏄ラ柡宓苯娈梺璺ㄥ櫐閿燂�????闂佹寧绻傛鍛婃櫠椤旂瓔娈介柣鎰皺婢ф稓绱掔紒妯肩畵闁崇粯鎹囧畷褰掝敊閻ｅ奔鎲鹃梻鍌欑劍鐎笛兠哄澶婄柧闁绘ǹ灏欓弳锔界節婵犲倻澧涢柡鍛箞閺屾稓浠﹂悙顒傛闂佹寧绋撻崰鏍涢崨鎼晝闁靛骏�????閿熺瓔妲遍梻浣告惈閻寰婇崜褏鐭夛�??锟姐儱鎳夐崼顏堟煕閺囨娅冪紒銊ヮ煼濮婃椽宕烽鈩冿�??锟介梺鎼炲妿婢ф寮查崼鏇熷殤妞ゆ帒鍊归敍蹇擃渻閵堝棙灏甸柛�?�枛�?�曟椽鏁愭径瀣幐闂佽法鍣﹂敓锟????闂佸摜濮甸悧鐘荤嵁閸愵喗鍊婚柦妯侯槺妤犲洤鈹戦悙鍙夘棞鐟滄壆鍋ら敓锟???妞ゅ繐妫涚壕浠嬫煕鐏炲墽鎳呴柛鏂跨У閵囧嫰濡搁妷褍鈪甸悗瑙勬磻閸楀啿顕ｉ敓�????????濠电姷鏁搁崑鐐哄垂閸洘鏅濋柍杞扮贰閻掍粙鏌嶉崫鍕舵�??閿熻姤绂嶅⿰鍫熺厵闁告繂瀚ˉ婊兠瑰⿰鍕姢妞ゎ亜鍟存俊鍫曞礃閵娿儱顫撳┑掳鍊楁慨鐢稿箖閸�?偛鏄ラ柣鎰惈缁狅綁鏌ㄩ弮鍥棄濞存粌缍婂娲礈閼碱剙甯ラ梺绋款儏閹冲氦顣鹃梺鍛婃处閸ㄩ亶鍩涢幋鐘电＜閻庯綆鍋掗崕銉╂煕鎼淬垹濮嶉柡宀嬬秮閸┾剝绻濋崒�???妗撻梻浣虹帛娓氭宕板Δ鍐╁床婵犻潧顑呯壕鍏肩�?婵犲倸顏柣锝囧厴濮婄粯鎷呴崨濠傛殘濠电偠顕滅粻鎾崇暦閹达箑�?嬫い鏍ㄧ☉閳ь剙鐏氶妵鍕箻閸楃偟浠鹃梺鎶芥敱閸ㄥ潡寮婚妶澶婄畳闁圭儤鍨垫竟鍕渻閵堝懐绠伴柣鎾愁煼�?�曞爼顢楁担鍝ユ濠电姰鍨奸崺鏍拷?锟介崶锟??�?夐柣鎴ｅГ閳锋垿鏌涘┑鍡楊�?鐞氼亪姊洪崨濠冪叆婵炴挳顥撻崚鎺撶節濮橆剛顦悷婊冾�?瀹曟垿骞樼紒妯轰画闂佸搫顦伴娆徫涘畝鍕拺闁告縿鍎辨牎濠电偛寮剁划鎾诲箠閻愮儤鐒硷�??锟姐儱妫�?▓銉╂⒑闂堟稓澧曢柛濠傛啞缁傚秵銈ｉ崘鈺冨幗闂佺粯鏌ㄩ幖顐︼�??锟芥總鍛婄厱闁绘柨鎼禒褏绱掓潏銊ョ闁归�???閺佹捇鏁撻敓�??????闂佺鍕垫當闁哄嫨鍎甸弻锝夊箛椤掍焦鍎撶紓浣哄�?�缂嶄線寮婚妸鈺佺睄闁搞儺鐓堝Λ鍕箾鐎涙鐭婄紓宥咃工椤繐煤椤忓嫭宓嶅銈嗘尵婵绮敓鐘崇厽闁靛繆鏅涢悘鈩冦亜閵娿儲鍤囬柛鈹垮灲楠炴ê煤缂佹ɑ娅嶉梻浣虹帛椤洭寮幖浣规櫖婵犲﹤瀚换鍡涙煏閸繄绠抽柛鎺嶅嵆閺屾盯鎮ゆ担鍝ヤ桓閻庢鍠栭崯鍧椼偑娴兼潙閱囬柣鏂挎惈楠炴劙姊绘担鍛婂暈濞撴碍顨婂畷鏉款潩椤戠偞妞介獮�???顢欓悾灞藉箞闂備礁鍟块幖顐﹀疮椤愶絿顩烽弶鍫厛濞堜粙鏌ｉ幇顒佲枙闁稿孩妫冮弻鈩冩媴缁嬪簱鍋撻崸�???绠板┑鐘插暙缁剁偤鏌涢埄鍐︿沪濠㈣娲樻穱濠囨�?��?�割喖鍓扮紓浣靛妼閻栫厧鐣烽幋锟??绠荤紓浣姑禒顓㈡⒑閸濆嫷妲规い鎴炵懃铻為敓�????閸曨兘鎷洪梺鍛婄缚閸庤鲸鐗庢俊鐐拷?锟介崝灞轿涘┑鍡╁殨闁哄被鍎卞敮闂侀潧顦崹娲棘閳ь剟姊绘担铏瑰笡闁挎岸鏌ｈ箛鏂垮摵鐎殿喗濞婇崺锟犲川椤�?儳骞堥梺璇插嚱缂嶅棝宕滃▎蹇�?瘎婵犵數鍋涢悺銊у垝鎼淬垻浠氶梻浣哥枃椤曆囨煀閿濆宓佹俊顖濇閺嗭箓鏌涢妷銏℃珔闁绘劕锕濠氬磼濞嗘埈妲梺鍦拡閸嬪棛鍒掗弮鍫濊摕闁靛鍎抽ˇ�???鏌ｆ惔顖滅У闁告挻鑹鹃悾鐑藉蓟閵夛妇鍘遍梺鏂ユ櫅閸熶即鍩婇弴銏＄厽闁规儳顕幊鍛磼鏉堛劍灏伴柟宄版嚇濡啫鈽夊顐ｅ亝闂傚�?�绀�?幖顐︻敄閸℃瑧鐭欓柟鍓х帛閸庡銇勮箛鎾跺缂佺姵姘ㄩ幉闈╂嫹?閿熺瓔鍠栫壕濠氭煏韫囧�????閿熶粙鎮″☉銏℃櫢闁跨噦�????闁诲函缍嗛崜娑溾叺濠德帮�??锟芥慨鐑藉磻濞戞◤娲敇閳ь兘鍋撴担鑲濇棃宕ㄩ鐙呯床婵犵數鍋為崹鍫曟偡閵夆晛鍑犳繛鎴炃氶弨浠嬫煟濡櫣浠涢柡鍡忔櫊閺屾冻�????閿熺瓔鍋嗗ú�?�橆殽閻愯宸ラ柣锝嗙箞瀹曠喖顢曢姀鈶╁亾椤撱垺鈷戦柤鎭掑剭椤忓煻鍥寠婢舵鍔烽梺鍝勭▉閸樹粙鎮￠敐澶屽彄闁搞儯鍔岄崵顒佺箾閸忕厧濮ч柟鍑ゆ�??闂佽法鍠曟慨銈吤洪弽顓勫洭鎮界粙鑳憰闂佸搫娲ㄩ崰鎾剁不妤ｅ啯鐓曟い顓熷灥閺嬫稑鈹戦鑺ョ婵﹨娅ｇ槐鎺懳熼懖鈺冪獥闂備焦鎮堕崝蹇撐涢崟顖ょ稏闊洦鎷嬪ú顏嶆晜闁告侗鍘洪悽濠氭⒒娴ｅ憡鎯堟い锔垮嵆閺佹捇鏁撻敓�???????闂傚倸鍊搁崐鐑芥嚄閸洖绠犻柟鎹愵嚙閸氬綊鏌″搴�?�箹缂佺媴锟?????婵犵數濮烽弫鍛婃叏閻戣棄鏋侀柛娑橈攻閸欏繘鏌熺紒銏犳灍闁稿骸顦…鍧楁嚋闂堟稑顫�?紓浣哄珡閸パ咁啇闁诲孩绋掕摫閻忓浚鍘奸湁婵犲﹤鎳庢禍鎯庨崶褝韬�?┑鈥崇埣瀹曠喖顢�?悙宸拷?锟介梻鍌欑閹诧繝鎮烽妷褎宕叉慨妞诲亾鐎殿喖顭烽弫鎰緞婵犲嫷鍚呴梻浣瑰缁诲�?�螞椤撶倣娑㈠礋椤撶姷锛滈梺璇�?��?�閸愶絾瀵栫紓鍌欑贰閸ｎ噣宕归幎钘夌闁靛繒濮Σ鍫ユ煏韫囨洖啸妞ゆ挻妞藉铏圭磼濡搫顫嶅銈嗘⒐閻楃姴顕ｉ幎鑺ユ櫢闁绘ê鍟块�?顒傛暬閹嘲鈻庤箛鎿冧痪缂備讲鍋撻柛鎰靛枟閻撶喖鏌熼崹顔碱伀缂佲檧鍋撻柣搴㈩問閸犳牠鈥﹂悜钘夌畺闁靛繈鍊曢敓�????????婵犵數濮烽�?�钘壩ｉ崨鏉戝�?�闂傚牊绋撻弳锕傛煟閵忊懚褰掓儗濡ゅ懏鐓曢柍鈺佸暟閳洟鏌嶉柨�?�伌闁哄瞼鍠栭幊鏍煛娴ｉ鎹曞┑鐘殿暜缁辨洟寮查銈嗩潟闁圭儤姊癸拷?锟芥岸鏌熺紒妯虹瑲婵炲牐顕ц灃闁绘﹢娼ф禒婊堟煟濡や焦灏板ǎ鍥э躬楠炴牗鎷呴懖婵勫妽閵囧嫰寮�?崶顭戞缂傚倸鍊归幑鍥ь潖缂佹ɑ濯撮柧蹇撶畭閳ь剙锕弻娑㈠箻鐎靛摜鐤勯梺闈涙閸熸潙鐣烽妸鈺婃晬婵犲ň鍋撶紒锟??顦甸幃妤冩喆閸曨剛顦ュ┑鐐茬湴閸斿孩绔熼弴銏″癄濠㈣绻傜紞濠囧极閹版澘鐐婇柍鍝勶拷?锟介崯鎺楁⒒娴ｈ鍋犻柛濠冪墵閹兘鏁傞悾灞告敵婵犵數濮村ù鍌炲极閸愵喗鐓ユ繝闈涙婢跺嫰鏌涢幒鎾舵创婵﹨娅ｉ崠鏍即閻斿憡绶梻浣呵归鍡涘箰閹间緤锟???閿熶粙宕�?鍢壯囨煕閳╁喚娈橀柣鐔稿姉缁辨挻鎷呯粵瀣櫍缂備胶绮换鍌炴偩閻戠瓔鏁嶆繝闈涚墢閺夌ǹ鈹戦悙鏉戠仸闁荤啙鍥у偍闂侇剙绉甸埛鎴犵磽娴ｇ櫢�????閿熶粙骞嬮敓�????�???鍫熸叏濮�?棗鍘撮柡瀣⒐缁绘繃绻濋崒婊冾杸闂佺粯鎸婚悷锕傚Φ閸曨垰妫�?悹鍥ㄥ絻椤牆鈹戦悙棰濆殝缂佺姵鎸搁悾鐑藉箣閿燂�??缁犳稒銇勯弮鍌涘殌濞存粓绠栭弻锝夋偄閸涘﹦鍑″銈冨劚缁绘﹢寮诲☉銏″亹闁归鐒﹂悾鑲╃磽娴ｆ垝鍚柛�?�仱楠炲棝寮崼鐔告珳闂佹悶鍎�?弲顏嗘閹惰姤鈷掑ù锝呮嚈瑜版帒�?�夋い鎺戝閸嬶紕鎲搁弬璺ㄦ殾婵犻潧妫崥�?�熆鐠轰警鍎忛柣婵囨濮婃椽宕ㄦ繝搴㈢暭闂佺ǹ顑嗛崝娆忣嚕閵娾晜鍤嶉柕澶涚导缁ㄥ姊洪崫鍕犻柛鏂块叄閸╁﹪寮撮�?鈽呮�??閿熶粙鐓崶銉ュ姢闁伙絿鏁婚弻鈥崇暆鐎ｎ剛锛熸繛瀵稿婵″洭骞忛悩瑁佺櫢�????閿熺瓔浜欐竟鏇炩攽閻樼粯娑фい鎴濇搐閻ｅ灚鎷呴幖鐐╁亾閹烘埈娼╅柨婵嗘噸婢规洘淇婇妶鍥ラ柛�?�仧閺侇噣鏁撻悩闈涚ウ闁诲函缍嗘禍鏍绩娴犲鐓曢柣锟??娼ч�?�濂告煕閵娿儳浠㈡い顐㈢箳缁辨帒螣閼测晜鍤岄梻渚婃嫹?閿熻棄鑻晶顔姐亜椤撶偞绌挎い锔界叀閹藉爼鎮欑紙鐘电畾闂�?潧鐗嗛幊蹇涘闯濞差亝鐓涢柛娑卞枤缁犳牠鏌曢崶褍顏紒鐘崇洴楠炴﹢骞囨担椋庣濠电姷鏁搁崑娑㈠触鐎ｎ喗鍋嬫俊銈呭暞瀹曞弶绻涢幋鐑囦緵闁哥喎鎳忛妵鍕籍閸パ冩優闂佺儵鏅涳拷?锟解晝鎹㈠☉姘棜閻庯綆浜欏Ч妤呮煥閻曞�?�锟????闂傚倷绀�?幖顐�?嫉閿燂拷?鐓ゆ俊顖欒閸ゆ鏌涢弴銊ョ仩闂佸崬娲︾换婵嬫濞戞瑯妫炲銈冨劜缁诲牆顫忕紒妯诲�?�闁荤喖鍋婇崵�?�磽娴ｇ瓔鍤欓柛濠呭劵濡喐绻涳拷?锟界ǹ甯堕柣掳鍔戝畷鎴�?磼閻愬鍘搁梺鎼炲劘閸庨亶鎮�?鍫熺厽闁规儳宕崝锕傛煛锟??瀣М鐎殿噯锟???????????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜忛弳锕傛煟閵忊懚鍦玻濡ゅ懏鐓曢柍鈺佸暟閳藉鐥幆褎鍋ラ柡宀嬬秮閿燂�??闁斥晛鍟禒鈺呮⒑闁偛鑻崢鍝ョ磼閳ь剚绗熼�?顒勬晲閻愭祴�?介悗锝庡亜濞堟繈姊洪崜鑼�?帥闁稿鎳橀幃鐢稿礃濞村锟??闂佺粯锕╅崰鏍倶鏉堛劎绠惧璺侯儑濞叉挳鏌℃担绋挎殻濠碉拷?锟界埣�?�曞爼鍩￠崘銊ь唽濠电姷鏁搁崑鐐哄垂閸洘鏅搁柨鐕傛嫹???闂傚倸鍊烽悞锕傛儑瑜版帒鍨傞柦妯侯樈閻掔晫鎲稿澶嬪仱妞ゆ挶鍨洪埛鎴︽偣閸ャ劌绲绘い鎺嬪灲閺屾盯骞嬪┑鍫⑿ㄩ悗瑙勬礃婵炲﹪寮幇顓炵窞濠电姴瀚弳鏉库攽閻愬瓨灏伴柛鈺佸暣�?�曟垿骞欓崟�???�????闂佽法鍠曟慨銈吤哄⿰鍫濆偍鐟滄棃宕洪悙鍝勭闁挎洍鍋撻敓�????閸愵喗鐓冮柛婵嗗閳ь剛鎳撻�?�鍧�?箣濠靛啯�???闂佹寧绋戯拷?锟筋剚绂嶆總鍛婄厱濠电姴鍟版晶顏呫亜椤愩垻绠洪柕鍥ㄥ姍楠炴帡骞嬪┑鍡橆吇缂傚倸鍊搁崐鐑芥倿閿曞偊�????閿熶粙宕堕浣镐画闁荤喐鐟ワ�??锟筋喚绮绘ィ鍐╃厵閻庢稒顭囬幊鍐煟韫囷絼閭柡�?嬬秮楠炴﹫锟???閿熻姤顭囬ˇ浼存⒑閸濆嫮鐏遍柛鐘崇墵閻涱噣宕卞鍏硷拷?锟介梻浣规偠閸婃宕伴幇顔藉床婵炴垯鍨圭粻鐢告煙閻戞ɑ鈷愰柟鎻掋偢濮婃椽妫冨☉娆愭倷闂佽法鍣﹂敓锟??????闂傚倷鐒︼拷?锟窖呯矙閹寸姭鍋撳鐓庡籍鐎规洝娅曪�??锟界》锟???閿熻姤锚閳ь剛鏁婚幃宄扳枎韫囨搩浠鹃梺璺ㄥ櫐閿燂拷??闂佽姘﹂～澶娒洪敃鍌氱闁绘梻鍘ч弰銉╂煏婢舵稓鐣辩紒鍓佸仜閳规垿鎮欓棃娑楀闂佽楠搁…鐑藉蓟閿濆牏锟??闁哄洨鍋樺▽顏堟⒑缁嬪灝顒㈠┑鐐诧躬閵嗕線寮�?崼婵囧祶濡炪倖鎸炬慨鐑芥晬濠靛鈷戠紒�?�锟??浼存煠瑜版帞鐣洪柛鈹惧亾濡炪倖甯婇悞锕傚磹閹邦喒鍋撶憴鍕闁告梹鐟╅獮鍐ㄢ堪閸喎�???????闂傚倸鍊烽悞锔兼�??閿熺獤鍥ㄦ櫢闁跨噦锟??????闂傚倷绀�?幖顐�?箯鐎ｎ偆顩叉い蹇撳濞兼牜绱撴担鑲℃垶鍒婏拷?锟藉摜纾兼繛鎴烇供閸庡繑绻涢崼顐㈠箻缂佽鲸鎸婚幏鍛存惞閻熸壆顐奸梻浣告啞濮婄懓煤閻旂厧绠栧Δ锝呭暞閸婅崵绱掑☉姗嗗剱闁哄懌鍨藉娲川婵犲啫顦╅梺绋款儏濡繂鐣烽�?銈呯妞ゆ棁袙閹疯櫣绱掔紒銏犲箹闁瑰啿绻�?弫鎾绘晸閿燂�??????闂佽法鍣﹂敓�?????闂佸憡娲﹂崑鍛存倵椤掍胶�???闁汇垽娼у瓭濠电偠顕滅粻鎾诲箖閿熺姴鍗抽柣鏃囨閻�?牓姊婚崒姘卞�?缂佸甯¤棢婵犲﹤瀚ㄦ禍婊堢叓閸パ屽劀闁瑰嚖锟???闂佽法鍠嶇划娆忣嚕婵犳碍鏅搁柨鐕傛嫹??闂佹寧绻傛鍛婄濠靛鍊堕煫鍥风到瀵噣鏌＄仦鐣屝ら柟鍙夋尦�?�曠喖顢曢妶鍕闂佽姘﹂～澶娒洪悢鍝ヮ洸闁割偅娲栭弰銉╂煃閳轰礁鏆炲┑顖涙尦閹綊宕堕柨瀣�??闂佽法鍠曟慨銈夊磻閹达附鈷掗柛灞捐壘閳ь剚鎮傚畷鎰槹鎼达絿鐒奸梺璺ㄥ櫐閿燂拷??濡ょ姷鍋為悧鐘伙�??锟介弴銏犖ч柛鈩冦仦缁剝淇婇悙顏庢嫹?閿熶粙宕濊缁骞嬮悩宸闂佺鍕垫當缂佺嫏鍥ㄧ厱妞ゆ劧绲块。鍙夌箾閸涱厽鎼愰柍钘夘�?楠炴ê鐣烽崶鍠插洦鐓涢敓锟???鐎ｎ剛袦闂佽鍠撻崹鑽ゅ垝濞嗘挸绠伴幖杈剧到濞村洭姊洪懡銈呮瀾缂侇喖瀛╅弲璺何旈崘鈺傛濠德帮拷?锟介幊搴ㄦ偪妤ｅ啯鐓涢悘鐐额嚙閸�?粓鏌ｉ幘瀛樼缂佺粯鐩獮�?�攽閸℃艾鐓橀梻浣告惈椤戞垶淇婇崶顒佸剦妞ゅ繐鐗滈弫鍥ㄧ箾閹寸伝鍏肩珶閺囥垺鈷掗柛灞捐壘閳ь剚鎮傚畷鎰槹鎼达絿鐒奸梺璺ㄥ櫐閿燂�???濡ょ姷鍋涢ˇ闈涱�?�闁�?秵鐓欑紒娑橆儏娴滅増鎱ㄦ繝鍛仩闁归锟??閸ㄩ箖鎼归銈勯偗闂傚�?�鑳舵灙闁挎洏鍎甸獮鍐磼閻愬瓨娅滈梺缁樺姇婢у酣鎮块�?�???鈹戦悙鏉戠仸闁荤噦绠撳畷鏇㈩敂閸啿鎷洪梻鍌氱墐閺呮盯鎯佸⿰鍫熺厱婵せ鍋撶紒鐘崇墵楠炲啴鏁撻悩鑼啋缂傚�?�鐒﹁彜闁归攱妞藉娲閳轰胶妲ｉ梺鍛娚戦崝娆忕暦閻戠瓔鏁囨繛鎴灻兼竟鏇炩攽閻愭潙鐏﹂悽顖涱殔閳诲秵绻濋崘鐐啍闂佺粯鍔樼亸娆戠不婵犳碍鐓涢悘鐐跺Г椤ユ粍銇勯幘鐐藉仮鐎规洝绮剧粻娑㈠棘濞嗗彞绱梻鍌氾�??锟介崐椋庣矆閿燂�??閺佹捇鏁撻敓�??????闂備浇顕э�??锟解晝绮欓崼銉ョ柧婵犲﹤鍠氶崵妤呮煕閺囥劌鐏犻敓�????鐎ｎ偁浜滈柡宥冨妿閵嗘帡鏌涢敓锟???娴滃爼寮婚敐鍡樺劅妞ゆ牗绮庢牎濠电偛鐡ㄧ划搴ㄥ礂閿燂�??閹繝顢楅崟鍨櫌闂佸憡娲﹂崜娑㈠储閽樺鏀介柣鎰綑閻忋儻�????閿熻姤娲﹂崜鐔奉嚕閹间焦鏅滈柛鎾�?拑绱查梻浣虹帛閿氱痪缁㈠弮閸┿儲寰勯幇顓犲帗闂佽姤锚椤﹁棄危閹间焦鐓冮悹鍥ㄧ�?閸欏嫭顨ラ悙鍙夊枠妞ゃ垺枪椤﹂亶鏌燂�??锟界ǹ鍘存慨濠傤煼瀹曟帒顫濋悙�???�????闂佽法鍠曞Λ鍕箒闂佹悶鍎滈埀顒勫几閺嶎厽鐓涢柛銉ｅ劚閻忊晠姊婚崒銈呯仸闁哄被鍔戝鎾�?�閸ャ劌�????闂佽法鍠撻弲顐ゅ垝婵犳凹鏁嶉柣鎰嚟閸欏棝姊虹紒妯荤闁稿﹤缍婇弫鎾绘晸閿燂�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崘鐐暥閻炴碍绻堝缁樻媴閸涘﹤鏆堥梺鍦�?归悥鐓庣暦濠靛绠ｉ柨锟??鍎崇粊锕傛椤愩垺澶勭紒瀣浮�?�煡骞栨担鍦�????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殘閳ь剙绠嶉崕鍗灻洪妶澶婂瀭婵犻潧娲ㄧ粻楣冩煕閳╁喚娈曠紒鍌氼儐缁绘盯宕楅懖鈺侇潷缂備胶绮粙鎴︻敊韫囨侗鏁婇柤濮愶拷?锟介崵顒勬⒒娴ｅ憡鎯堥柟鍐茬箻楠炲啴宕掗悙鑼舵憰闂侀潧艌閺呮粓宕戦崱娑欑厱閻忕偛澧介埥澶愭煥閻曞倹锟????缂傚倸鍊搁崐鎼佸磹閹间礁纾瑰�?�捣閻棝鏌ㄩ悤鍌涘?闁芥ɑ绻堝娲敆閳ь剛绮旈幘顔煎嚑濞撴埃鍋撻柟顔肩秺�?�曞爼顢旈崟顓燁嚄闂備礁鎼Λ瀵哥不閹捐钃熼柨鐔哄Т閻愬﹪鏌嶆潪鎵妽闁诲氦宕电槐鎾存媴缁嬫鏆㈤梺绋款儍閸婃繈鐛�?崘銊庢棃宕ㄩ鑺ョ彸闂備礁鎲￠崝鎴﹀礉锟??鍕舵�??閿熶粙宕卞▎鎴狅紳婵炶揪缍佸褎淇婇崗绗轰簻妞ゆ挾鍋涘Σ濠氭懚閻愮儤鐓曟繛鎴炵懄閸庢鏌℃担绋挎殻闁哄矉锟??????婵＄偑鍊ч懙褰掑疾閻樺樊娼栨繛宸簼閸嬶繝鏌ｉ敓锟???閻楀﹪宕伴幇鐗堚拺缂佸顑欓崕鎰版煙閻熺増鎼愭い鏇秮閹崇娀顢楁担鍝ワ紡闂佽崵鍋炵粙鍫ュ礈濠靛缍栵�??锟姐儱顦伴埛鎴︽⒒閸喓娲撮柣娑欑矌缁辨帗娼忛妸锔绢槹閻庤娲忛崹铏圭矉閹烘柡鍋撻敐搴�?�簮闁归攱妞藉娲閳轰胶妲ｉ梺鍛娒妶绋跨暦濠靛牃鍋撻敐搴�?�簽缂佺�?绠栭弻娑樷枎韫囷絾楔婵犫拃灞藉缂佽鲸甯″畷鎺戭潩濮ｆ瑣鍎甸弻鏇㈠炊閵娿儱顫掑Δ鐘靛仦鐢繝鐛Ο鍏煎磯闁告繂�?�悷鏌ユ⒒娴ｈ棄鍚归柛鐘冲姉閸掓帒顓奸崶褍鐏婇梺瑙勫劤绾绢參寮抽敂鐣岀瘈濠电姴鍊搁弳濠囨煛鐎ｎ亪鍙勯柡�???鍠撻�?顒傛暩鏋亸蹇曠磽娴ｈ娈旀い锔炬暬楠炲啫螖閸涱垰绁﹂梺鍓茬厛閸犳牗鎱ㄦ惔鈽嗘富闁靛牆绻愰惁婊堟煕閵娿劍鐝紒鏃傚枛瀵挳锟??閻樼粯鏆呮繝寰峰府锟???閿熶粙鎳楅崼鏇炲偍闁告鍋愰弨浠嬪箳閹惰棄纾归柡鍥ュ灩閻ゎ喗銇勯幇鍓佺暠闁绘帒鐏氶妵鍕箳閹搭垰濮涢梺鍛婂笂閸楁娊寮诲澶嬪癄濠㈣埖蓱绗戦梺鍙ョ串缂嶄礁顫忓ú顏勫瀭妞ゆ洖鎳庨崜鎶芥⒑闁偛鑻晶顔姐亜椤撶偛妲婚摶鐐烘煕濞戞瑦鍎楅柡浣稿暣閺屾洝绠涙繝鍌氣拤闂佽鍠楅悷鈺侇潖濞差亜绠伴幖娣�?灮閿涙﹢姊虹粙鎸庢崳闁轰礁顭烽悰�???宕橀妸搴嫹?闂佺粯鎸堕崐鏍Φ閸曨喚锟??闁圭偓娼欏▍婵嬫⒑瑜版帗鏁辨俊鐐舵椤繑绻濆顒傦紲濠殿喗锚�?�曨剟路閳ь剛绱撻崒娆戭槮妞ゆ垵妫濋獮鎰板礈瑜嶉崹婵嗏攽閻樺磭顣查柛濠勫厴閺岋綁骞嬮悜鍡欏姺闂佸憡枪妞村摜鎹㈠┑�?�仺闂傚牊�???閵忋倖鐓曢柣鏂挎惈椤ｅジ鏌￠崨顓犲煟闁诡喕绮欏畷銊︾�?閸曨偄绠為梻鍌欑閸熷潡骞栭锟??纾归悹鍥梿閾忓厜鍋撳☉娆欎緵婵炲牅绮欓弻锝夊箛椤掍讲鏋欓梺绋垮濡啴寮婚埄鍐╁�?�闂傚牃鏅滈敓锟????闂佽法鍠嶇划娆撶嵁閸愵喖�?堢憸灞解柦椤忓牊鐓㈡俊顖欒濡叉椽鏌ｉ妶鍛仾缂佺粯绻堥幃浠嬫濞磋翰鍎甸弻鈩冩媴閸涘﹤鏆堢紓浣虹帛閻╊垶宕洪埀顒併亜閹哄秷鍏岀紒鐘冲劤闇夐柨婵嗘噹閺嗛亶鏌涘顒碱亪鍩ユ径濞㈢喎饪伴崟顒夋閻庤娲︽禍婵嬪箯閸涱垱鍠嗛柛鏇ㄥ墰瑜板棝姊婚崒姘炬嫹?閿熺晫绮堥敓�????瀹曨垶宕搁敓�????缁犺銇勯幇鍓佺暠缂佺姷�???閻擃偊宕堕妸褉濮囬梺绋款儏閸婂潡寮诲☉銏犵疀闁稿繐鎽滈崙褰掓⒑閸濄儱校闁告梹鐗滈幑銏犫攽閸モ晝鐦堥梺绋挎湰缁矂銆傞敓锟?????闂備礁澹婇崑鍡涘窗閹惧墎涓嶅Δ锝呭暞閻撴洟鏌嶉埡浣稿絹闁瑰濮抽悞濠偯归悡搴ｆ憼闁绘挻娲熼幃妤呮晲鎼存繃鍠氶梺璺ㄥ櫐閿燂拷??闂傚倷绀�?幖顐︽儗婢跺瞼绀婂�?�姘ｅ亾闁绘侗鍣ｉ弫鎾绘晸閿燂拷??闂佸湱鍘х紞濠囷拷?锟介弴銏℃櫜闁告稑鐡ㄩ敍妤呮⒒閸屾熬�????閿熺晫绮堥敓�????楠炴牠顢曢埗鑺ョ〒閳ь剟娼ч幗婊勭▔瀹ュ鐓欓柟瑙勫姦閸ゆ瑩鏌﹂崘顏勬灈闁哄矉缍佸顒勫垂椤�?枻锟???閿熶粙姊虹粙娆惧剰妞ゆ垵顦靛璇测槈閵忊晜鏅濋梺闈涚墕閹冲繘鎮橀敓锟???濮婃椽宕ㄦ繝鍌滃帎缂備胶绮换鍌烇綖韫囨稒鎯為悷娆忓绾绢垶姊洪棃娴ㄥ綊宕曢弻銉�?仧闁靛繈鍊栭埛鎴︽煟閻斿憡绶叉繛鍫�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾剧懓顪冿拷?锟筋亝鎹ｉ柣顓炴闇夐柨婵嗘噺鐠愶繝鏌ｅ┑濠冪�?�闁宠鍨块幃鈺呭矗婢跺⿴妲遍梻浣呵归鍛村磹閸ф钃熸繛鎴欏焺閺佸啴鏌ｅΟ璇茬祷濠殿喖娴风槐鎺楁�?�閿燂拷?閸斻倖銇勯鐘插幋鐎殿喛顕ч埥澶愬閻樻彃绁梻锟??娼ф灙闁稿氦娅曪拷?锟藉ジ宕堕浣叉嫼闁哄鍋炴竟鍡浰囬敃鍌涚厱濠电姴鍊归崑銉�??閿熺瓔鍠栭�?�閿嬩繆閹间礁鐓涢柛灞剧煯缁ㄤ粙姊绘担鍛靛綊寮甸鍕櫢闁跨噦锟???????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归崷顓犱笉閻犲洩顥嗚ぐ鎺撴櫜闁割偒鍋呯紞鍫ユ⒑闂堟稒澶勭紒璇插暣婵＄敻宕熼姘兼綂闂佹枼鏅涢崰姘涢崘顔斤�??锟介悷娆忓绾炬悂鏌涢敓�????閸ㄥ潡濡存担鑲濈喓鎮伴埄鍐╂澑闂備礁澹婇崑鍡涘窗閹邦儷鎺撴償閵婏腹鎷婚梺绋挎湰閻旑剟骞忛敓锟????闂佽法鍠嶇划娆忕暦閹邦収妲归幖杈剧悼閿燂�????婵°�?�濮烽崑鐐烘偋閻樹紮�????閿熶粙寮村杈┬㈤梻浣规偠閸庢椽宕滃▎鎴犱笉闁靛�?璐熸禍婊堟煛閸愵煉锟???閿熶粙宕甸埀顒佺箾鐎涙鐭婂褏鏅Σ鎰板箳閹宠櫕姊归幏鍛偘閳╁喚娼旈梻鍌欒兌鏋柨鏇橈�??锟介垾锟??鐣￠柇锟??娈ㄦ繛鏉戝悑濞兼瑧澹曟總鍛婄厽闁归偊鍠涜棢闂佺懓鍢查…宄邦潖閾忓湱鐭欓柟绋垮閹烽亶姊洪悡搴ｇШ缂佺姵鐗犻弫鎾绘晸閿燂�???婵＄偑鍊栫敮鎺楀磹閹间礁鍌ㄩ柟缁㈠枟閻撴瑦銇勯敓�????閸庤櫕绂掗柆宥嗙厸濞达絿枪閺嗭綇�????閿熻姤娲樼敮鎺楋綖濠靛洦缍囬柍鍝勶拷?锟介惁鎺楁⒒閸屾熬锟???閿熺晫绮堟担鍦彾濠电姴娲ょ壕濠氭煕濞戝崬濮告繛宸簻閿燂拷?濡炪倖鎸鹃崑娑㈡倵椤撱垺鈷戠紒�?�锟??鐗堛亜閺囶澀鎲撅�??锟筋噮鍣ｅ畷濂告偄閸涘﹦褰囨繝鐢靛仦閹稿鎳濇ィ鍐╂櫇妞ゅ繐鐗婇崑妯荤節婵犲倸顏紒鐘荤畺閹鈽夊▎妯煎姺闂佹椿鍘奸敃锔炬閹炬剚鍚嬮柛婊冨暢閸氼偊鎮�?▓鍨灕妞ゆ泦鍥х�?濠㈣埖鍔曢～鍛存煟濡吋鏆╅柡澶嬫�?�濮婂宕掑顑藉亾閹间焦鍋嬪┑鐘插閻瑩鏌熼悜姗嗘畷闁稿﹤澧庨埀�???绠嶉崕閬嵥囨导鏉戠厱闁瑰濮风壕濂告倵閿濆骸浜介柛搴涘劦閺屾稒鎯旈敍鍕姱闂佸搫鐭夌换婵嗙暦閵娾晩鏁婇柣鎰靛墮閿燂拷?????婵犳鍠栭敃銉ヮ渻娴犲宓侀柟閭�?幗閸庣喖鏌ㄥ┑鍡樺窛闁哄棎鍊濆缁樻媴閻戞ê娈岄梺鍝ュ枎濞硷繝寮绘繝鍥ㄦ櫜闁告粈绀佸▓銊╂⒑鐟欏嫬鍔跺┑顔猴拷?锟藉畷鎴�?礋椤栨稓鍘遍棅顐㈡处閼圭偓绂嶈ぐ鎺撶厱婵☆垰�?遍惌娆愭叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚�?�鑳舵灙闁挎洏鍊濋獮澶愭晬閸曨厾鐒块悗骞垮劚椤︻垳绮诲杈ㄥ枑濠㈣埖鍔曠紒鈺伱归悩宸剱闁绘挾鍠愭穱濠囶敍濠靛浂浠╂繛�?�稿У閻╊垶寮婚敓鐘插耿闊洦姊归悵姘舵煥閻曞倹锟???????闂佽法鍣﹂敓�??????闂佽法鍣﹂敓�?????????闂備礁鎼ú銊╁磻閻旇櫣鐭撻柣姘摠閿燂拷??闂佽法鍠曟慨銈吤洪弽顓炍х紒�?�儥閸ゆ洟鏌熺紒銏犳灍闁稿�?�伴弻褍顫濋敓锟???閳ь剙顭峰顐ｃ偅閸愨斁鎷婚梺绋挎湰閻熝囧礉�?�ュ鍊电紒妤佺☉閸樻儳煤椤忓嫬鍞ㄥ銈嗘尵閸嬬喖鏁嶅▎鎾粹拺闁告稑锕︾紓姘舵煕鎼淬劋鎲鹃挊鐔告叏濡灝鐓愰柣鎾寸懅缁辨帪锟???閿熺瓔鍘界涵鍫曟煛閸曨偓�????閿熶粙婀佸┑鐘诧工鐎氼噣鎯岄幒妤佺厽闁瑰灝鍟禍甯�??閿熻姤娲栭悥鍏间繆閹间焦鏅搁柨鐕傛嫹?闂傚倸顦粔鐟邦潖濞差亝顥堥柍鍝勫暙閸╁矂姊虹涵鍛撶紒顔奸鍗遍柟鐗堟緲缁犳娊鏌ㄩ悤鍌涘?闁诲孩纰嶅畝鎼佸蓟濞戞ǚ鏋庨煫鍥风稻閳绘挸鈹戦埥鍡椾壕缂佺姵鎸搁～蹇撁洪鍕炊闂佸憡娲﹂崜姘跺箯閸楃偐鏀介柣鎰硾閻ㄦ椽鏌涢悩鏌ュ弰闁诡噣绠栭幃婊堟嚍閵夈儰绨甸梺鍦帶閻°劏鎽梺璺ㄥ櫐閿燂�???闂傚倸鍊风粈浣圭珶婵犲洤纾诲〒姘ｅ亾鐎规洘妞藉畷鐔碱敍濮樺啿鐓樻繝鐢靛仜濡﹥绂嶅┑瀣厱闁圭儤鍤氳ぐ鎺撴櫜闁告侗鍠栭弳鍫ユ⒑閸濄儱鏋旈柛�?��??锟介獮鍐╃鐎ｅ灚鏅�?┑顔缴戝畷锟??宕ラ锔斤拷?锟介悷娆忓缁岃法绱掔紒妯肩疄闁绘侗鍠楅幆鏃堝Ω閿燂拷?閻у嫭绻濋�?锝嗙【閻庢稈鏅犻獮澶愭偋閸垻鐦堥梺姹囧灲濞佳勭閿曞�?�鐓曟い顓熷灥閻忥讣�????閿熻姤娲滈幊鎾跺弲濡炪�?�绻愶拷?锟筋噣鏁嶅☉銏♀拺缂侇垱娲栨晶鍙夈亜閿曞倻绱伴柕鍥ㄥ姍楠炴帡骞橈�??锟芥褰搁梻鍌欑閹测剝绗熷Δ鍛獥婵°倕鎳庣粣妤呮煙闁箑骞樼紒鐘荤畺閹鎮介惂鏄忣潐閻�?酣姊绘担绛嬪殐闁哥姵鐗犲畷鎰板锤濡ゅ啫绁﹂梺鍛婂姂閸擃噣寮崼婵堝姦濡炪倖甯掞拷?锟筋剟鎮″┑瀣厵闁硅鍔﹂崵娆撴煕閵娿儻锟???閿熶粙濡甸崟顖氱睄闁稿本绋掗悵顏呯箾鐎涙鐭婇柣鏍帶椤繒绱掑Ο璇诧�??锟介梺鎯х箳閹虫挾绮敓鐘斥拺闁荤喓澧楅崯鐐烘煙閸涘﹤鈻曪�??锟芥洩锟???濠碉紕鍋戦崐鏍ь啅婵犳艾纾婚柟鎯у濡垳绱撴担闈涚仼鐎殿噮鍠氶�?顒侇問閸犳绻涙繝鍥ф瀬闁稿本绋掗崣蹇涙煙闁缚绨介柣鈺侀叄濮婄粯鎷呯粵�?�秷濠电姰鍨鸿摫闁哄懓鍩栭幆鏃堝Ω閿燂拷?娴犲ジ姊绘笟鍥у缂佸鎸抽幊婊呮喆閸曗晙绨婚梺鍝勭▉閸嬪嫭绂掗敃鍌涚厱閻庯�?�鍐ㄢ拤缂備胶绮换鍐崲濠靛纾兼慨姗嗗幗椤斿秶绱撻崒娆掑厡濠殿喗鎸抽垾锕傛�?�閽樺鎽曢梺鏂ユ櫅閸燁垱鍒婇幘顔界厱婵犻潧瀚崜楣冩煏韫囧﹥顫婃繛鍫㈠閵囧嫯绠涢幘铏閻庤鎸稿Λ鎾箯閿燂�???闂佽法鍠曟慨銈吤洪弽顓炍ч柟闂寸缁犳牠鏌曡箛瀣舵�??閿熶粙鎯岄敓�????椤法鎹勭悰锛勬箙婵炴潙鍚嬮悧鐘差潖婵犳艾纾兼慨妯煎亾閿燂拷??闂佽法鍠撻弲顐ゅ垝閸儲鏅搁柨鐕傛嫹?濡ょ姷鍋涢ˇ鐢稿极瀹ュ绀嬫い鎾跺Х閸橆垶姊绘担渚敯闁规椿浜浠嬪礋椤栨氨鏌у┑鐘绘涧椤戝棝鎮￠妷鈺傛櫢闁跨噦�????????缂傚倸鍊烽懗鑸垫叏閻戣姤鏅搁柨鐕傛嫹?闂備礁鎼張顒勬儎椤栫偟宓侀柛銉墮鎯熼梺鎸庢婵倗娆㈤鐐╂�?闁绘劘灏欓幗鐘电磼椤旇偐肖闁告帗甯￠獮妯兼嫚閼艰埖鎲伴梻�???娼ц墝闁哄懏绋撻悮鎯ь吋婢跺鍘遍梺闈涱槶閸斿秶娑甸悙顒傜闁割偒鍋勫顔芥叏婵犲懏顏犻柟椋庡█閹崇�?顢楅崒婊勬緰闂傚倷鑳舵灙婵炲鍏樺顐ゆ嫚�?�割喖娈ㄩ柣鐘叉搐濡﹪宕ワ�??锟筋亶鐔嗛柤鍝ョ仚閹达箑鐤炬繝濠傜墛閳锋垹绱掗娑欑濠�?勭叀閺岋綁鎮㈤弶鎴斿亾濠靛绠归柣鐔煎亰閸熷懏鎱ㄦ繝鍐噰婵﹤顭峰畷鎺戭潩閻愵剙锟???闂佽法鍠嶇划娆忕暦閹版澘绠瑰ù锝呮憸閿涙瑩姊鸿ぐ鎺擄紵閿燂�??娴ｅ搫顥氱憸鐗堝笚閻撴瑩姊婚崒姘煎殶妞わ讣濡囬惀顏堝箚瑜忕粔娲煛閿燂拷?閸犳牕顫忛懡銈傚亾闂堟稑顥忔俊宸枤缁辨帡鎮欓敓�????閸斻倗绱撳鍜冭含鐎殿喖顭烽幃銏ゅ礂鐏忔牗�?�介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閿燂�???闂佹寧绻傛鍛婃櫠娴煎瓨鐓熼柨鏇�?亾闁绘鎹囬獮鍐ㄎ旈崘鈺佹�?�闂佸憡娲﹂崜娑⑺囬妷鈺傗拺缂備焦顭囨晶顏堟煕濮橆剦鍎愮紒宀冮哺缁绘繈宕堕妸銉㈠亾婵犳碍鐓㈡俊顖滃皑缁辨岸鏌曟繛褍�?�弸鎴︽煥閻曞倹锟???闂佸憡娲﹂崑鍡涙偩濞差亝鈷戦柟绋挎捣缁犳挻绻涚仦鍌氬濠㈣娲樼粋鎺炴嫹?閿熺瓔鍋嗛崢閬嶆煟韫囨洖浠滃褌绮欓獮濠囧幢濡晲绨婚梺鍝勶�??锟介娆徫熼�?顒勬煥閻曞�?�锟???????婵＄偑鍊栭崝褏寰婇悾灞筋棜闁规儼濮ら埛鎴︽煕濠靛棗顏敓�????娴煎瓨鐓熼柍鍝勶工閻忥箓鏌曢崱鏇犵獢鐎殿喗鎸抽敓�????闁斥晛鍟悵鎶芥⒒娴ｈ鍋犻柛搴㈢矌娴狅箓骞嗚閻忓酣姊婚崒姘炬�??閿熶粙宕愰悜鑺ユ櫢闁跨噦�???????闂傚倷鑳舵灙妞ゆ垵妫濋獮鎰板箹娴ｅ湱鐣抽梻鍌欒兌缁垶鏁嬪┑鈽嗗灠閿曨亜鐣烽弴銏犵疀闁绘鐗忛崢浠嬫⒑鐟欏嫬鍔ら柣掳鍔庣划鍫嫹?閿熺瓔鍠楅悡娆愩亜閿燂拷?閺嬪鎳撻崸妤佺厵妞ゆ梻鏅幊鍥殽閻愬瓨宕屾鐐村浮�?�曞崬螣閾忚楔濠电姷鏁告慨鐢割敊閺嶎厼绐楁俊銈呭缂嶆﹢姊绘担鍛婂暈闁哄被鍔戦弻濠囨晲婢跺苯绁︽繝銏ｅ煐閸�?洜绮婚悷鎳婂綊鏁愰崶銊ユ畬婵炲瓨绮撴禍璺侯潖濞差亜绀堥柟缁樺笂缁ㄨ偐绱撴担绛嬪殭閻庢矮鍗抽獮鍐倻閽樺鎽曢梺闈涱檧閼靛綊骞忛搹鍦＝濞达絽澹婇崕蹇涙煟韫囨梻绠炴い銏☆殜閿燂拷?閹鸿櫕绂嶅⿰鍫熺厪濠电偛鐏濋崝婊勩亜閵壯冧户缂佽鲸甯掗悾婵嬪礃椤斿吋鎳欑紓鍌欒兌缁垳鎹㈤崼婵堟殾闁割偅娲嶉�?顒佺墵椤㈡牠顢楅�?�???煤閿曞�?�鍋傞柡鍥ュ灪閸婂爼鏌ｉ幇顓炵祷闁抽攱妫冮弻锝夊箼閸愩劎浠╁銈庡弨濞夋洟骞夐幘顔肩妞ゆ帒鍋嗗Σ鏉库攽閻戝洨鍒版繛灞傦拷?锟介弫鍐敂閸繄鐣哄┑鐐叉閹尖晠寮崒鐐寸厱闁哄洦锚婵＄厧霉濠婂牏鐣洪柡灞炬礋�?�曠厧鈹戦崶鑸碉骏婵＄偑鍊愰弲娑橆嚕閸撲焦宕叉繝闈涙川閿燂拷?闂佺ǹ鏈划宀勶拷?锟藉ú顏呪拺婵懓娲ら�?顑撅�??锟藉畷浼村冀椤撶喓鐣抽梻鍌欒兌鏋紒缁樺姍�?�曘儻锟???閿熺瓔鍓涚粈濠囨煙鏉堥箖妾柣鎾跺枛閺岀喖鎮滃Ο铏逛患婵炲濮甸惄顖炲蓟閺囥垹鐐婄憸宥夘敂椤撶噥娈介柣鎰綑濞搭喗顨ラ悙宸剶妞ゃ垺绋戦～婵嬵敆婢跺绁紓鍌氾拷?锟介崐鎼佸磹妞嬪海鐭嗗�?�姘ｅ亾閽樻繈姊婚崼鐔剁繁闁绘帞鏅幉鎼佸棘閸栤槄锟???閿熻棄霉閿濆洨銆婇敓�????娴犲鐓熸俊顖涱儥閸ゅ�????閿熻姤鎮堕崕鐢稿箖閿燂拷?椤繈鎮℃惔銏㈠綆闂備浇顕栭崹浼存儗閸岀偟宓�?柟鐑樺殾閿燂�??閹峰懘宕崟顐ゎ吋婵犵绱曢崑鎴�?磹閺嶎厽鍋嬫俊銈呮噺閸嬶紕鎲歌箛鏇炲灊闁挎繂顦Λ�???骞栵�??锟芥ɑ灏伴柡鍌�?亾闂傚�?�鐒﹂弸濂稿疾濞戙垹鐤い鏍仜绾惧綊鏌熼幍顔碱暭闁绘挻娲熼弻宥夊传閸曢潧鍓抽梺璺ㄥ櫐閿燂拷??闂佽姘﹂～澶娒洪敓�????閺佹捇鏁撻敓�??????闂傚倷绀�?幉锟犲礉閹达箑绀夐幖鎼厛閺佸﹪鏌涢妷顔煎闁抽攱甯￠弻娑氫沪閹规劕�????闂佺粯鍨兼慨銈夊吹閸曨垱鐓曢柟鎹愬皺閸斿秹鏌涜箛鏃傜煉闁哄本鐩、鏇㈡晲閸℃瑯妲梺璺ㄥ櫐閿燂拷??闂佸壊鍋嗛崰鎾跺姬閳ь剟姊婚崒姘卞�?濞撴碍顨婂畷鏇炵暆閸曨剛鍘撻悷婊勭矒瀹曟粓濡歌娑撳秹鏌熼幆褏锛嶉柡鍡畵閺屾盯顢曢敐鍡楊槱闂佽桨绀佸Λ妤呮箒闂佹寧绻傚В銉ф喆閸曨厾褰鹃梺鍦劋椤ㄥ棝鍩涢幒鎳ㄥ綊鏁愰崨顔兼殘闁荤姵鍔х换婵嬪蓟濞戞瑦鍎熸繛鎴ｆ珪閿燂�???闂佽法鍠嶇划娆愪繆閹绢喖�?冩い鏃傚帶閼板灝鈹戦悙鏉戠仸闁荤喆鍎茬粋宥呂旈埀顒勫煘閹达附鍊烽柡澶嬪灩娴犙囨⒑閹肩偛濡芥俊鐐舵椤曪綁寮婚妷銉ь啇婵炶揪绲藉﹢閬嶅矗閸℃稒鈷戠紓浣股戦敓�????闂佽法鍣﹂敓�????????闂傚倸鍊搁崐鎼佸磹妞嬪孩顐芥慨妯挎硾閻掑灚銇勯幒鎴�??閿熻姤绂掑⿰鍫熺厾婵炶尪顕ч悘锟犳煛閸涢偊鍟囬柟鍑ゆ嫹?闂佽法鍠撻弲顐ゆ兜閸洖纾婚柟鎹愬煐閸犲棝鏌涢弴銊ュ闁挎稒鐩娲川婵犲孩鐣锋繝鐢靛仜閿曨亪骞冩导�?�樻櫢闁跨噦�????闂佽法鍣﹂敓�???????闂佽法鍣﹂敓�?????闂佺ǹ鏈粙蹇旂濠婂牊鐓欓柟浣冩珪濞呭懘鏌ｈ箛锝勯偗闁哄本鐩幃鈺冪驳绾應鍋撻崸妤佺厸閿燂�??閳ь剟宕伴弽顓ㄦ嫹?閿熻棄鈻庨幘婢勨晠鏌曟径娑㈡闁诡喗鐟╁缁樻媴缁嬭儻鍩炲┑鐐叉▕閸欏啫顕ｆ繝姘櫜濠㈣泛锕ラˉ婵嬫⒑閸撹尙鍘涢柛鐘炽仦缁ㄧ儤绻濋悽闈浶ユい锝勭矙瀹曟粌鈹戦崶鈺冾啎婵犵數濮撮崑鍡楊焽閺嶎偆纾藉ù锝堝亗閹寸偛鍨旈柟缁㈠枟閻撴洘绻濋棃娑欘棞妞ゅ景鍛＝闁稿本绋掑畷灞炬叏婵犲懏顏犵紒顔界懇瀹曠ǹ螖閳ь剙顕ｉ悧鍫㈢閻庢稒顭囬惌搴㈢箾婢跺娲撮柟�???绠栭幃婊呯驳鐎ｎ偅娅栨繝鐢靛Т閿曘倧锟???閿熺瓔鍓涙竟鏇㈩敍閻愮补鎷洪梻鍌氱墛娑撶懓鈽夐姀鐘碉紲濠电姴锕ら幊蹇涘窗閹烘鈷掗柛灞捐壘閳ь剛鍏�?幃鐐烘晜閸忕厧锟???闂佽法鍠撻悰銈夊川椤旂厧绨ラ梻浣呵归惉濂稿磹濞戙垹鐐婇柕濞垮労閸ゃ�?�姊洪崫鍕垫Ч闁搞劌缍婂畷銏ゆ焼�?�ュ棌鎷洪梺闈╁瘜閸樺ジ宕濓�??锟筋喗鐓曢柕鍫濇娴溿垽鏌曢崶銊ュ妤犵偞甯￠獮姗堟�??閿熻姤顭囪ぐ鎼佹⒒閸屾瑧顦﹀鐟帮躬瀹曟垿宕ㄩ姘亰闂佽鍎煎Λ鍕不閼姐�?�纾藉ù锝堫嚃閻掍粙鏌涘鍡曢偗婵﹨娅ｉ崠鏍即閻愭祴鎷ゆ俊鐐�??锟介崝宀勫箠濡警鍤曢柟鎯板Г閺呮彃顭跨捄渚剳闁告﹫�?????闂佽鍑界紞鍡涘礈濞戞壕鍙烘繝寰峰府�????閿熻姤鎱ㄩ悜钘夌；闁绘劕鐏氶弳婊堟煥閻斿搫孝缂佺姵鐗楃换娑㈠幢濡闉嶉梺绋款儍閸旀垿寮诲☉顫�??閿熶粙骞嬪┑鍛嚬婵＄偑鍊栧褰掑箰閹间礁鐓�?柟�?�稿仜缁犵娀姊虹粙鍖℃敾妞ゃ劌妫濋獮鍫ュΩ閳哄偊锟???閿熶粙鏌�?Ο渚Ш闁挎稒鐩铏圭磼濡搫顫岄梺鍦拡閸嬪﹤鐣疯ぐ鎺戠＜闁绘劕顕崢鍗烆渻閵堝骸骞楅柛銊ф暬瀵悂濡舵径瀣幐闂佺硶妲呴崢楣冩偩閻㈠憡鐓涢敓�????閳ь剟宕伴弽顓ㄦ嫹?閿熻棄鈽夐姀鈽呮�??閿熶粙妫呴顐㈠箹闁哄鐗婄换婵堝枈婢跺锟???闂佽法鍠曞Λ鍕舵嫹?閿熻棄閰ｉ弻娑㈠籍閳ь剟宕归悽闈╃稏闊洦鎷嬪ú顏嶆晜闁告洦鍙庨崯鍥⒒娴ｈ櫣甯涢柛�???鐗滅划濠囧箻椤旇偐锛涢梺瑙勫礃椤曆囧礃閳ь剙顪冮妶搴�?�⒕闁瑰嚖锟???闂佽法鍠曟慨銈夊箚閸喆浜滄い鎰剁悼閻帡鏌ㄩ悤鍌涘�??婵＄偑鍊栫敮濠傤渻閹烘梹宕查柛鈩冪⊕閻撶喖鏌曡箛濠冨殙闁革富鍘鹃惌鍡涙�?�閿濆骸浜栧ù婊勭矒閺岋拷?锟筋吋閸愩劌顬夐梺姹囧妽閸ㄥ爼濡甸崟顖氭闁告煭銈呮儓婵犳鍠栭敃銉ヮ渻娴犲绠栭柣鎴ｆ缁犮儲銇勯弮鍥撻柛鐘崇墱缁辨捇宕掑▎鎰偘濡炪�?�娉﹂崨顖滅厠闂佹眹鍨婚弫鎼佹儗婢舵劖鐓欓柣鎴炆戠亸鐢告⒒閸曨偄顏柡灞剧☉閳藉顫滈崼婵嗩潬闂備礁鎲￠敃銏＄鐠轰警娼栨繛宸簼椤ュ牊绻涢幋锝夊摵妞ゅ骸妫濆濠氬磼濮橆剦浠奸柣搴㈠嚬閸犳绮嬪澶婄濞达綀顫夊▍鍡涙⒑閸忛棿鑸柛搴�?�船椤曪綁骞愭惔锝囩槇闂佹眹鍨藉褍鐡梻浣烘嚀閸熻法鎹㈤敓�????閵嗕線寮�?崼鐔蜂汗缂傚倷鐒﹂�?�鍥�?储闁�?秵鈷戦柛婵嗗琚梺鍛婃煥鐎涒晠寮查敓锟???????婵＄偑鍊栧Λ浣规叏閵堝洣鐒婇柨鏇烇�??锟介悡娆愩亜閺冨倹娅曢柟鍐插暣閺佹捇鏁撻敓锟???????婵＄偑鍊栭崝鎴﹀垂閺勫繈浜归柟顖ゆ嫹?�???浠嬫煟濡椿鍟忛柡鍡樼矌缁辨帗娼忛妸锔绢槹閻庤娲橀崹鍧楃嵁鐎ｎ喗鏅搁柨鐕傛�??缂佺偓鍎崇紞濠囧蓟閿燂拷????闂佽法鍣﹂敓�?????????闂備緤锟???閿熻棄鑻晶鎾煥閻曞�?�锟???婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划濠氬蓟閵夛妇鍘棅顐㈡搐椤戞垿骞忛敓�?????闂佽法鍠撻弲顐ゅ垝婵犳碍鏅查柛鈩冨姃缁ㄥ姊洪崫鍕犻柛鏂块叄閸┿儲寰勶�??锟姐劋锟??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏妞ゆ洝绮鹃ˇ褰掓煛閿燂拷?閸犳牕顫忛懡銈咁棜閻庯綆浜滅敮顖炴煟鎼淬値娼愰柟鍝ュ厴閹偤鏁傞悾灞告敵婵犵數濮村ù鍌炲极瀹ュ棛锟??闂傚牊绋掗ˉ娆愭叏鐟欏嫷娈樼紒杈ㄥ浮閹瑩顢楅�?顒勫礉閵堝鐓曟慨姗嗗墻閸庢劗绱掑畝鍐摵缂佺粯绻堝畷鍫曟嚋閸偅鐝梻鍌欒兌缁垶宕濋弴銏″仱闁靛ň鏅涘Ч鏌ユ煟濡偐甯涢柣鎾跺枛楠炴牠骞栭鐔虹獢婵炲瓨鍤庨崹鐑樼┍婵犲浂鏁冮柕蹇曞娴煎啴姊虹化鏇熸珖闁稿鍊濋悰顕嗘�??閿熺瓔鍠楅敓�????????闂傚倸鍊风粈�???宕ワ�??锟筋喖绠栭柛灞惧嚬閻掔晫鎲稿澶婄叀濠㈣泛�?�掑Ο鍕攽椤旂�?�榫氭繛鍜冪秮楠炴垿宕熼姣尖晠鏌曟径娑橆洭鐟滅増宀稿缁樻媴閻戞ê娈岄梺鎼烇�??锟介悧鐘荤嵁閿燂�????婵犵數濮烽弫鍛婃叏閻戣棄鏋侀柛娑橈攻閸欏繘鏌ｉ姀鐘差棌闁轰礁锕弻鈥愁吋鎼达�??锟界缂備焦鍔栭〃濠囧蓟閻旂厧绠查柟浼存涧濞堫厾绱掗悙锟??�?冩い顐㈩槹缁岃鲸绻濋崶顬囨煕鐏炲墽鐓瑙勬礋濮婄粯鎷呴崫銉︼�??锟藉┑鈽嗗亜鐎氭媽妫熼梺姹囧灮鏋紒鐘崇墵閺岋綁鏁愰崨顖�?紘闂佹椿鍘介悷鈺呭蓟濞戞粠妲煎銈冨妼閹虫ê顕ｉ銉ｄ汗闁圭儤鎸撮幏缁樼箾鏉堝墽鍒伴柟璇х節楠炲棝宕奸悢铏诡啎闁诲繒鍋涢崐鍛婃叏閸屾壕鍋撶憴鍕；闁告濞婇悰顔嘉熼崗鐓庣彴闂佸湱绮敮鎺撶閸洘鈷掗柛灞剧懅鐠愪即鏌涢幘瀵告噮缂侇喗妫冮幃鐣�?矙鐠恒劌骞堥梻浣烘嚀椤曨厽鎱ㄦ搴☆棜闁芥ê顥㈣ぐ鎺撴櫜闁告侗鍨抽弳娑㈡⒑闁偛鑻晶顖炴偨椤栥�?�锟??妤犵偛鍟撮幃婊堟寠婢跺矈鍚嬮梺璺ㄥ櫐閿燂�???????闂傚倸鍊搁崐椋庣矆閿燂拷?楠炴牠顢曢埛姘そ婵℃悂鍩℃担鐚寸幢闂備胶绮濠氬储瑜嶆晥闁哄被鍎查悡銉╂煛閸モ晛鍓抽柟鍑ゆ嫹?闂佽法鍠嶇划娆撳箖閿熺姴唯闁冲搫鍊婚崢浠嬫⒑閸濆嫭宸濋柛瀣舵�????????闂傚倸鍊搁崐鎼佸磹妞嬪孩顐芥慨妯挎硾閻掑灚銇勯幒鎴�??閿熻姤绂掑⿰鍫熺厾婵炶尪顕ч悘锟犳煛閸涱厾鍩ｏ�??锟芥洩绲惧鍕醇濠婂懐娉垮┑锛勫亼閸婃牠宕濋幋�???鏄ラ柛鏇拷?锟介敐澶婄濞达絿鎳撴禍妤呮⒑闂堟稓澧曟い锔垮嵆閹繝宕�?鐣屽幈濠电�?娼уΛ妤咁敂閳哄懏鏅搁柨鐕傛�??????闂備礁鎼ú銊╁磻濞戞氨妫憸蹇曟閹烘梻纾兼俊顖濆亹閻ゅ嫬鈹戦埥鍡椾簻闁哥噥鍋婇崺銉�?緞閹邦剛顢呴梺缁樺姈瑜板啴藟閹扮増鈷戦悹鍥у级閸炲銇勯銏╂█妤犵偞鍔栭ˇ鐗堟償閵忊晛浠烘繝娈垮枟閿氬褍楠搁悾鍨瑹閳ь剟寮婚垾鎰佸悑閹艰揪绲肩划鎾绘煙閸忓吋鍎楅柣鎾崇墦瀵偊宕卞☉娆戝帗閻熸粍绮撳畷婊冾潩椤撶姭鏀虫繝鐢靛Т閸熶即銆呴悜鑺ワ�??锟介柨婵嗛�?�娴滅偤鏌涢敓锟???娴滆泛顫忓ú顏咁棃婵炴垶鑹鹃�?�娲⒑绾懏鐝柛�???鐗犲鏌ュΨ閳哄�?�鎷绘繛杈剧到閹诧繝骞嗛崼銉︾厸闁割偒鍋勬晶�???鎮￠妶鍡曠箚妞ゆ牗鐟ㄩ鐔兼煕閵堝棭娈滈柡灞剧洴瀵挳濡搁妷銈囩埍婵犵鍓濊ぐ鍐偋閹捐钃熼柡鍥风磿閿燂拷?婵犵數濮撮崰姘焽閹达附鏅搁柨鐕傛嫹????缂傚倷绀�?ˇ閬嶅箠閹句紮缍栭煫鍥ㄧ⊕閹偤鏌涢敂璇插箻闁挎稒绮岄埞鎴�?煡閸℃浠撮梺绋款儐閸旀瑩骞冩ィ鍐╋�??锟芥俊顖濆亹閻﹀牓姊哄Ч鍥х伈婵炰匠鍕浄婵犲﹤鐗婇悡銉╂煛閸ヮ煉鍏柟鍑ゆ�??闂佽法鍠嶇划娆撳极閹扮増鍊烽柛鎾茶兌閺夋悂姊洪崫鍕窛濠殿喚鍏橀弫宥呪堪閸愶絾锟??闂佸疇妫勫Λ妤呮�?�閵夆晜鐓曢悗锝庡亜婵秹鏌熼娆戠獢鐎规洖銈告俊鐑芥晜閹冪闂傚倷绀�?崥�?�矈閹绢喖鐤鹃柣鎰煐閿涘倿姊婚崒娆戠瓘闁瑰嚖�????闂佽法鍠曞Λ鍕嚐椤栨稒娅犻柡灞诲劜閸婂爼鐓崶銊︹拻闁瑰啿娲弻鐔碱敍濮橆剦浠鹃梺璇″灡濡啯鎱ㄩ埀顒勬煏韫囧鐏俊鎻掓喘濮婄粯鎷呴崷顓熻弴闂佹悶鍔忓Λ鍕�??锟介崶顏嶆Ъ缂備礁鍊圭敮锟犲春閿熺姴纾兼俊顖氭贡閻╁酣姊绘担鍛婃儓婵炲眰鍔戝畷浼村箻缂佹ê鍓归梺璺ㄥ櫐閿燂拷??缂備浇椴哥敮锟狅�??锟藉▎鎴濇�?�閺夊牃鏅涢幃鎴炰繆閵堝洤啸闁稿鍋ら弫鍐閵堝洤绁﹂梺鎼炲劘閸斿秵鍒婇幘顔界厱婵炴垶菤閻鏌涘顓犳噭缂佺粯绻堥幃浠嬫濞磋翰鍎甸弻鈩冩媴閸涘﹤鏆堥梺閫涚┒閸�?垿骞冩禒瀣窛濠电姴鍊归悿鍕⒒娴ｈ櫣甯涢柛鏃撶畵�?�曟粌鈻庨幘宕囶槷闂佸搫鍟悧濠囧煕閹烘鐓曢悘鐐插⒔閹冲懏銇勯敂鑲╃暤闁哄本鐩幃銏ゆ煥鐎ｎ亙娣俊銈囧Х閸嬬偤鎮ч悩浼欐�??閿熶粙寮撮姀鈩冩珕闂佸吋浜介崕鏌ユ偟閺嶎厽鈷掑�?�姘ｅ亾婵炰匠鍥佸洭顢曢敓锟???閻ょ偓绻涢幋娆忕仾闁稿浜弻锝夊箛闂堟稑顫梺璺ㄥ櫐閿燂拷??婵犵數濮烽弫鍛婃叏閹绢喖纾圭紓浣股戝▍鐘崇箾閹存瑥鐏柣鎾冲暣濮婃椽宕归鍛壈闂佽绻戦幐鎶藉蓟閿涘嫪娌柛鎾�?嫬鍨辨俊銈囧Х閸嬬偤鏁冮姀�???鍤曢柛顐ｆ礀缁狅綁鏌ｅΟ鐓庝化闁稿鍓濈换婵嬫偨闂堟稐绮堕梺�?�︽澘濡块柛鎺撳笒椤撳ジ宕堕妸銉ョ哎闂備礁鎲￠崝锔界濠靛棛鏆﹂柛娆忣槺缁犻箖鏌燂拷?锟芥鎳冮柣蹇婃櫊閺岋綁顢橀悤浣圭暥濡炪値鍘煎锟犲箠濠婂牊鍋ㄦ繛鍫ｆ硶娴煎洭姊婚敓�????閳ь剛鍋涢懟顖涙櫠椤旂晫绠剧痪顓㈩棑閿燂拷?閻庢鍠涢褔鍩ユ径鎰潊闁绘﹢娼ч獮鎰版⒒娴ｅ懙褰掑嫉椤掑�?�鍨濓拷?锟姐儱顦粈鍡樼箾閹寸儐鐒搁柡鍐ㄧ墛閸嬫劙姊婚崼鐔衡棩缂侇喛娉涢—鍐Χ閸℃浠村銈忕畵濞佳囶敋閿濆鏁冮柨鏇楀亾缁炬儳銈搁弻锝夊箛椤撶喓绋囬梺璋庡啫顏紒缁樼箞閿燂拷?闁挎繂妫涢妴鎰版煥閻曞�?�锟???????闂備礁鎼悮顐﹀磿閺屻儱鐓曢柟鐑橆殕閻撴洟鎮�?悙鎻掆挃闁瑰啿�?�槐鎺撴媴閸濆嫷鏆梺闈涙搐鐎氭澘顕ｉ幘顔藉亜闁告繂�?�ч幏浼存煟鎼淬�?�娼愭繛鎻掔箻�?�曡绂掞拷?锟筋亞鐣洪梺鍛婃寙閸屾稑濯伴梻浣虹帛閸旓箓宕滃棰濇晩闁搞儺鍓氶埛鎺懨归敐鍛暈閻犳劧绻濋弻娑欐償濞戞ǚ鍋撳┑瀣祦闁归偊鍙庡Σ褰掑箹濞ｎ剙鐏╅幖鏉戯躬濮婅櫣鍖栭弴鐐测拤闂�?潧娲﹂惄顖氼嚕閵婏妇顩烽悗锝庡亞閸橀亶鏌ｈ箛鏇炰粶濠�?傜矙閵嗗倿寮婚妷锔惧幈闂佺粯鏌ㄩ幖顐ｇ闁秵鐓涢敓�????鐎ｎ剛袦濡ょ姷鍋為敃顐﹀箯閿燂拷??闂佽法鍠曞Λ鍕箟閿熺姴绀嗘繛鎴欏灪閳锋垿鎮归崶锝傚亾閾忣偆浜舵俊鐐�??锟介崝宀勬晝椤忓嫷鍤曟い鎰剁畱缁犳稒銇勯幘璺烘�?�闁告柨鎳樺娲�?�閽樺濮ら柣蹇撶箲閻熲晠骞嗛崟顒佸劅闁靛⿵鑵归幏缁樼箾鏉堝墽鎮奸柣鈩冩�?�曢潧鈻庨幋鐘碉紲缂傚�?�鐒﹂敋闁诲繐鐡ㄩ�?�銉╂�?�閺夋垵顫掑Δ鐘靛仜闁帮綁骞愭繝鍐ㄧ窞閹兼番鍨洪崯娲⒒閸屾瑨鍏岄柛�?�ㄥ姂�?�曟洘娼忛埡渚囨濡炪�?�鎸堕崹鐟靶ч弻銉︾厱闁斥晛鍟伴埊鏇㈡煕婵犲嫭鏆柡灞诲妼閳规垿宕卞☉鎵佸亾閿燂拷?椤儻顦遍柛妤佸▕�?�濡搁妷銏☆潔濠殿喗锕╅崜姘舵�?�閸績�?芥い鏃傦�??锟介弨缁樹繆閻愭壆鐭欙拷?锟筋喖顭峰畷顭掓�??閿熻姤锚閳ь剛鍏橀弻銈夋嚌閻楀牏銆愬銈呮禋閸樼晫鎹㈠┑�?�櫢闁跨噦�????闂佸憡鍔戦崝澶愬箰閸愵亞纾藉ù锝勭矙閸濇椽鏌熼崨濠冿拷?锟芥い銏∩戠缓鐣�?矙閸喚鐛╂俊鐐拷?锟藉ú鏍箠韫囨稒鏅ù锝堟绾句粙鏌涚仦鍓ф噮妞わ讣�??????缂傚倸鍊风粈�???藝闁�?秴绠犻柟鍓х帛閸嬧晠姊洪崹顕呭剳闂傚嫬瀚槐鎺炴嫹?閿熺瓔浜炴禒顫�??閿熻姤鎸稿Λ婵嗩潖閾忓湱纾兼俊顖涙た濮婂灝鈹戦悙�?�樺碍閿燂拷?闁秵鍤嶉梺�???绉甸崑銊╂煕濞戞☉鍫ュ箯缂佹绠鹃弶鍫濆⒔閸掍即鏌熼搹顐ゆ噰鐎规洜鍏�?、锟??鎮㈠畡鎵搸闂佽法鍣﹂敓�????????闂備胶绮幐璇裁洪悢鐓庤摕婵炴垯鍩勯弫鍐煥濠靛棙鎼愭い鈺婂墴濮婃椽宕崟闈涘壉闂佸搫琚崝鎴濓耿閿燂拷?濮婅櫣绱掑Ο蹇ｄ簻铻ｅ┑鐘叉搐绾惧潡鏌熼幍顔碱暭闁绘挾鍠栭弻鐔煎箲閹邦厾銆愰梺鍝勵儐閻╊垶寮婚敓鐘虫櫢闁跨噦锟???闂佸摜濮甸悧鐘差嚕婵犳艾鐐婃い鎺嶇劍濞呭洭姊洪柅鐐茶嫰婢ф挳鏌熼鏂わ�??锟介柟顔规櫇缁辨帒螣閻撳骸绠洪梻鍌欑窔濞佳勭仚闂佸憡鏌ㄧ粔褰掞拷?锟介弮鍫熷亹闁汇垻鏁搁敍婊堟煛婢跺﹦澧戦柛鏂胯嫰闇夋い鏇�?亾闁哄瞼鍠栭、娆戞喆閸曨剛褰呮俊鐐�??锟介弻銊ф崲閿燂拷?閵嗕礁鈻庨幘宕囩暰閻熸粌閰ｅ畷鎰邦敍閻愮补鎷婚梺绋挎湰閻熝囁囬敃鍌涚厵缁炬澘宕禍浼存煙椤栨凹妲圭紒铏规櫕缁瑧鎹勯妸褍鐐婇梻鍌欑閹碱偆绮欓敓�????瀹曘垼銇愰幒鎴犲姦濡炪�?�鍨煎▔鏇⑺囬敃鍌涚厓閻犲洦鐓￠崣鍕殽閻愯揪鑰匡拷?锟筋喖鐖奸獮瀣堪閸曨偂绨奸梻鍌欐祰椤曆勵殽閹间礁鍌ㄦ繝濠傜墕绾惧鏌熼崜褏甯涢柣鎾冲暟閹茬ǹ饪伴崼婵堫槶闂佺粯姊婚崢褏绮婚弽顓熺厓闁宠桨�?�?弳娆戠磼閸撲礁浠遍柡�???鍠栭弻鍥晝閳ь剟鐛幇鐗堢厵闂佸灝顑嗛妵婵囨叏婵犲啯銇濋柟绛圭節婵�?�爼宕ㄩ閿亾閻愵剛锟??闁靛繈鍨洪敓�????濠碘槅鍋呯换鍫濐嚕椤愩埄鍚嬮柛锟??�?�?幃鎴炵節閵忥絾纭炬い鎴濇喘�?�曘垽鏌嗗鍡欏幗闁瑰吋鎯岄崹宕囩矈閻戣姤鐓曢柡鍌濇硶閻掓悂鏌ㄩ悤鍌涘?婵＄偑鍊栫敮濠囨嚄閼稿灚娅犳い鎺戯拷?锟界壕纭锋嫹?閿熻В鍋撻柛鎰靛枛閹界數绱撴担铏瑰笡缂佽鐗嗛悾鐑藉醇閺囩倣鈺呮煏婢跺牆鐏╁ù婊勫劤閳规垿鎮╁畷鍥舵殹闂佺粯鎸鹃敓锟???闁哄瞼鍠栭�?�锟??鎮㈡搴ｆ噯闂備礁鎲″鍦垝�?�ュ洦宕叉繛鎴欏灩�?�告繃銇勯幘璺烘珡婵☆偁鍊楃槐鎾存媴娴犲鎽甸梺鍦归�?�鐑界嵁韫囨稑宸濋柡澶嬪灦�?�撳秴顪冮妶鍡樺鞍缂佸甯￠敐鐐差吋閸℃洜绠氶梺缁樺姦娴滅兘骞忛敓锟????闂佽法鍠嶇划娆忕暦閿燂拷?????濠电偛顕崢褔顢氶銏℃櫢闁跨噦�???????婵＄偑鍊栧Λ浣肝涢敓锟????婵犵數濮电喊宥夋偂閻樼粯鐓欐い鎾跺枎缁楁帡鏌涢敓�????椤ㄥ﹪寮婚悢椋庢殝闂侇叏濡囬崥�?�攽椤旂�?�榫氭繛鍜冪悼閸掓帒鈻庨幘宕囶唶闁瑰吋鐣崹鐚存�??閿熻姤濞婂缁樻媴閾忕懓绗�?�┑鈽嗗亜缁绘ê鐣峰⿰鍫熷亜闁兼祴鏅涚粊锕傛椤愩垺澶勭紒瀣浮�?�煡骞栨担鍦�????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖骞戦幇闈涙闂佹眹鍊楅崑鎾诲Φ閸曨垰绠涢柍鍝勵儐閿燂�???闂佽法鍠嶇划娆忕暦閻熸壋�?介悗锝庡亞閸樺崬顪冮妶鍡�?濠殿喗鎸冲畷婵嗏堪閸喓鍘搁梺鍛婁緱閸犳宕愰幇鐗堢厸閻忕偠顕ф慨鍌炴煙椤旂尨锟???閿熻棄鐣烽幒鎴旀婵妫旈敓锟????婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙盯姊虹紒妯哄闁稿簺鍊濆畷鎴嫹?閿熺瓔鍠楅悡鐔镐繆椤栨繂鍚归敓锟???娴犲鐓冪憸婊堝礂濞戞碍顐芥慨姗嗗墻閸ゆ洟鏌熺紒銏犳灈妞ゎ偄鎳橀弻宥夊煛娴ｅ憡娈插銈呯箳閸犳牕顫忕紒妯诲�?�闁兼亽鍎抽妴濠囨⒑闂堚晝绉剁紒鐘虫崌閺佹捇鏁撻敓锟???????缂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛顐ｆ礀绾惧鏌熼幑鎰靛殭缁炬崘娉曢�?顒冾潐濞叉牕煤閵娧呯焼濠电姴鍊甸弨浠嬫煟濡搫绾ч柟鍏煎姍閺岋箓宕�?鍕拷?锟界紓浣虹帛閻╊垶鐛拷?锟筋亖鏋庨煫鍥ㄦ�?婵爼姊绘担鑺ワ�??锟介敓锟???閿燂�??瀹曨垶骞�?鑹版憰闂侀潧枪閸庮噣寮ㄦ禒瀣厱闁斥晛鍠涙笟娑欎繆椤愮媴锟???閿熶粙鈥旈崘顔嘉ч煫鍥ㄦ皑椤︿即姊虹粙鍧楋�??锟界痪缁㈠幖鍗遍柟鐗堟緲缁犺櫕淇婇妶鍕瓘闁瑰嚖�????闂佽法鍠曟慨銈夊Φ閸曨垰绠抽柛鈩冦仦婢规洟姊绘担鍛婂暈闁哄矉缍佸畷鎰旈崘鈺婃綗闂佸湱鍋撻崜姘跺触鐎ｎ喗鐓曟繝濠傚暙閺嗐垽鏌涘鐓庝喊闁诡喗顨呴埢鎾诲垂椤旂晫浜俊鐐拷?锟介崢楣冨礂濡櫣鏆﹂悷娆忓閸嬪懘鏌涢幇鈺佸闁汇倐鍋撴繝鐢靛仩閹活亞寰婃禒�?�疅闁跨喓濮寸壕瑙勩亜閺嶎偄浠﹂柍閿嬪笒闇夐柨婵嗘噺閸熺偤鏌涢悢鍝勪粶闁靛棙甯掗～婵嬵敇瑜庨悿�???鎮楃憴鍕缂傚秴锕妴浣糕槈濡嘲鐗氶梺鍛婂姂閸斿孩绂嶆导瀛樷拻濞达絽�?卞﹢浠嬫煕閵娿儳绉烘鐐差樀閺佹捇鎮╅崘韫暗闂備胶绮濠氬储瑜忕划鑽ゆ喆閸曨厾顔曢梺鎸庣箓妤犲憡鏅堕敓锟???閺岋�?绠涢敐鍛彎闂佸搫鏈惄顖炲箖閵忋�?�浼犻柕澶堝劚缂佲晠姊绘担鍛婃儓閻炴凹鍋婂畷婵嬪箣閿燂拷?缁犳牠鏌曢崼婵愭Ц缁炬儳鍚嬬换娑㈠箣閻戝洣绶甸梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煁妞ゃ劊鍎甸幃娆欐嫹?閿熺晫枪閳綊鏌ら幐搴�?�闁靛洤�?�伴獮鎺�?幢濡炴儳顥氭繝鐢靛Х椤ｎ噣骞忛敓锟????闂佽法鍠庨～鏇㈠磻閵忋�?�鐓涢敓�????鐎ｎ剛袦濡ょ姷鍋炵敮锟犵嵁鐎ｎ喗鍋愰弶鍫氭櫊閳瑰繘姊婚崒娆戠獢婵炰匠鍏犳椽濡惰箛鏂款�??闂佽法鍠愰崹婵嬪�?閹惰姤鍋樻い鏇楀亾妤犵偞甯￠弫鎾绘晸閿燂�???缂備胶濯寸徊鍓ф崲濠靛顥堟繛鎴炆戝▓顓熺箾鐎涙鐭婂褏鏅Σ鎰板箳閻愭潙�????闂佽法鍠撻悺�???绂嶉悙宸僵闁靛ň鏅滈悡娑㈡�?�閿濆簼绨介弫鍫ユ⒑缂佹ɑ鎯勯柛�?�工閻ｇ兘宕奸弴鐐嶁晠鏌ㄩ弮鍥舵綈閻庢氨鏅槐鎾诲磼濞嗘帒鍘￠梺璺ㄥ櫐閿燂�???缂傚倷鑳舵慨鐢告偋閻樺樊鍤曢悹鍥ㄧゴ濡插牊绻濇繝鍌涘櫧闁哄鎮傚娲传閸曨剙绐涢梺绋款儐缁嬫帞绮嬮幒鎳崇喖鎳￠妶鍥╂婵犵數鍋涢悧鍡涙倶濠靛鍑犳繛鎴炵懀娴滄粓鏌ㄩ弴姘樂闁告凹鍋呮穱濠囧矗婢跺﹤顫掑Δ鐘靛仦鐢繝鐛Ο灏栧亾闂堟稒鎲搁懖鏍⒒閸屾瑧绐旀繛浣冲嫮浠氶梻浣呵癸�??锟解晜绻涙繝鍥锋�??閿熶粙寮介鐐碉紲闂佺粯鍔楃悰銉╁箯濞差亝鈷掑�?�姘搐娴滅偤鏌涳拷?锟筋偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備礁鎲￠幐鍡涘川椤栥�?�闂梺璇查缁犲秹宕曢柆宥呯疇闊洦铔嬫径鎰�??锟介柣銏㈡暩閿涙粓姊虹粙鎸庢拱婵ǜ鍔忛崐鎾⒒娴ｅ憡璐￠柟铏尵閳ь剚鍑归崣鍐嵁韫囨稑宸濋柡澶嬪灥�?�撳棝姊虹紒妯忣亜顕ｉ崼鏇燂�??锟介柛顐犲劜閳锋垹绱掗娑欑闁哄缍婇弻娑虫嫹?閿熺瓔鍋呯亸顓熴亜椤忓嫬鏆ｅ┑鈥崇埣瀹曞崬螖閸愵亝鍣梻浣筋嚙鐎涒晠宕欒ぐ鎺戠煑闁告劦鍠栭弰銉︾箾閹存瑥鐏╃紒鐙呯秮閺岋絽螣閸忓吋姣勯梺鎸庣⊕缁矂鈥旈崘顔嘉ч柛鈩冪懃椤呯磽娴ｅ壊鍎愰悽顖滃仧閸掓帡宕奸妷銉ь槰濡炪倖姊婚弲顐﹀储閸涘﹦�???闁靛骏绲剧涵楣冩煥閺囶亜顩紒顔芥煥鐓ゆい蹇撴噽閸樻悂鏌ｈ箛鏇炰粶濠�?傜矙婵℃挳骞掑Δ浣哄帗閻熸粍绮撳畷婊堝Ω瑜忕粈濠囨煕閳╁啰鈽夌痪鎯ь煼閺屾稑鈽夐崡鐐典户闂佺粯甯掗敃銉╁Φ閸曨垰绠婚悹铏瑰劋閻庮厽绻涳拷?锟芥鐭嬬紒顔肩Ч婵＄敻宕熼鍓ф澑闂佸湱鍋撻崜姘婵傚憡鈷戦柛婵嗗閿涙梻绱掗煫顓犵煓闁糕晝鍋ら獮�?�晝閳ь剟鎮樺畷鍥ｅ亾鐟欏嫭�???婵炲眰鍊濋幃锟犳偄閸忕�?�锟???閿熶粙鎮峰▎蹇擃仾閿燂拷?閳ь剟鎮楃憴鍕�?闁告挻绻堥幃锟??宕橀瑙ｆ嫼闂佸憡绋戦敃銈嗘叏閿燂拷?闇夋繝濠傚缁犵儑锟???閿熻姤娲樻繛濠囷�??锟藉☉銏★拷?锟界紒顔款潐鐎氳棄鈹戦悙鑸靛涧缂佹彃娼￠幃娲籍閸繂鎯炲┑鐐叉閹稿宕愰崹顐ょ闁瑰鍋涚粭姘箾閸涱厸搴烽柟鍑ゆ嫹?闂佽法鍠曟慨銈吤洪敓�????閹兘濡搁埡浣勶箓鏌熼悧鍫熺凡缂佺姵濞婇弻鐕傛嫹?閿熺晫枪鍟搁梺鍛婏供閸撶喎顫忕紒妯诲闁告稑锕ら弳鍫ユ⒑閸涘﹥顥栫紒鐘虫尭閻ｉ攱瀵奸弶鎴濆敤濡炪倖鍔戦崐鎾剁箔婢舵劖鈷戦柛婵嗗閳诲鏌涘Ο鍦煓闁诡噯绻濇俊鐑藉煛閸屾粌骞楅梻浣告惈閸婄櫢锟???閿熺獤鍥х畾闁割偒鍓氶敓锟????闂佽法鍠曟慨銈囨崲閸儱钃熸繛鎴欏灪閸婂鏌涢埄鍐炬畼濞寸姷枪閳规垿顢欑涵閿嬫暰濠碉紕鍋犲Λ鍕偩閻戣姤鏅搁柨鐕傛�??閻庤娲╃徊鎯ь嚗閸曨厸鍋撻敐搴濈盎濠㈢懓绉瑰濠氬磼濞嗘帒鍘￠柡瀣典邯閺屻劑寮村Ο琛�?�亾濠靛鐏抽柨鏇楀亾闁伙綇绻濋獮宥夘敊閼恒儺鍟庨梻鍌欑窔濞佳勵殽韫囨洘顫曢柡鍥ｅ亾閳ь剙鎳橀幃婊堟嚍閵夈儮鍋撻悽鍛婄叆婵犻潧妫濋锟??霉濠婂嫬濮嶉柡锟??鍠栭弻顭掓嫹?閿熺瓔鍋佹禒銏犫攽椤旂�?�鏀绘俊鐐舵閻ｇ兘濡搁敂鍓х槇闂佸憡娲﹂崢楣冨汲閵堝鈷戦悹鍥ㄥ絻椤掋垻鐥弶璺ㄐф鐐插暣�?�曟帡鎮欓棃娑氥偊闂傚⿴鍋勫ú锔剧矙閹烘鐤鹃柟闂寸劍閿燂�?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖鎮ч崼鐔哄嚒闂佸憡鍨规慨鎾煘閹达附鍋愰悗鍦Т椤ユ繄绱撴担鍝勶拷?锟介柛銊ョ埣瀵濡搁埡鍌氫簽闂佺ǹ鏈粙鎴︻敂閿燂拷??闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖宕滆鐢盯鏌涳拷?锟筋偓鑰块柡灞炬礋�?�曠厧鈹戦幇顓夛箓姊虹紒妯哄闁挎洩绠撻獮澶婎潰閿燂�??閿燂�??濠电偞鍨舵灙闁硅姤娲熷娲礈閹绘帊绨撮梺绋垮閻擄繝宕哄☉銏犵闁绘鏁搁敍婵囩箾鏉堝墽鍒版い顐ｇ墵椤㈡棃宕ㄩ鐓庝紟濠电姰鍨奸崺鏍礉閺嶎厽鍋傞柡鍥ュ灩缁犲綊鎮�?☉娆樼劷闁宠棄顦甸弻宥堫檨闁告挻姘ㄩ幑銏ゅ醇閵壯冪ウ闂佸憡鍔﹂崰妤呭疾閹间焦鐓熸俊顖氭惈閺嗗崬霉濠婂嫮鐭掓慨濠冩そ�?�曟鎳栭埞鍨沪闂備礁鎼幊蹇曠矙閺嶎厼桅闁圭増婢樼粈瀣亜閺嶃劎鈻撻柟閿嬫そ濮婅櫣娑甸崨顓濇睏闂佺ǹ顑嗛惄顖氱暦濠靛鏅滃┑顔藉姃缁ㄥ姊洪棃娑辨闂傚嫬瀚悾宄扮暆鐎ｎ偄锟???闂佽法鍠曟慨銈吤哄Ο铏规殕闁归棿绀佺粻鏍喐閺傝法鏆﹀┑鍌溓归～鍛存煏韫囧﹥娅呴柡鍜佸弮濮婂宕掑▎鎴М闂佽绁撮崜婵堢箔閻旇偤鏃堝川椤撶偛浜堕梻浣虹帛閸旓箓宕滃顑芥�?�闊洦绋掗埛鎺楁煕鐏炲墽鎳呮い锔肩畵閺�?喓鍠婇崡鐐扮凹閻庡灚婢橈�??锟芥澘鐣烽崼鏇熸櫢闁跨噦�????闂佺粯甯掗悘姘跺Φ閸曨垰绠抽柛鈩冦仦婢规洜绱撴担绋库挃闁惧繐閰ｅ畷锝夊礃椤垵娈ㄩ梺瑙勫劶濡嫰鐛�?�?锛勭闁瑰鍋熼幊鍛存煕濡粯宕岄柟顔煎槻楗即宕熼鐘靛帨闁诲氦顫夊ú妯煎垝閹捐绠栭柕蹇婃濡插綊骞栧ǎ�???鐏い锟??娲熷缁樻媴閾忕懓绗″銈冨妼閹虫﹢骞冭缁绘繈宕惰閿涚喖姊虹紒妯荤叆闁告艾顑夐幃陇绠涢幘顖涙杸闂佺粯枪鐏忔瑧绮婚幎鑺ョ厽闁挎繂鎳庨懜褰掓婢舵劖鐓熸俊顖濇�???鎾煕鐎ｃ劌鐏柟渚垮妽缁绘繈宕ㄩ鍛摋闂備礁�?遍幊鎿勬�??閿熺晫澧楁穱濠囧箹娴ｈ�?�銊╂煥閺傚灝缍栫紒銊ョ摠缁绘繈鎮介棃娴讹絾銇勯敓锟???閻楃姴鐣锋导鏉戝唨妞ゆ挆鍕珨婵＄偑鍊栭幐鍫曞垂濞差亜纾垮璺侯儍娴滄粓鐓崶銊�?鞍缂佷讲鏅滄穱濠囶敍濮橆剦浼冨┑顔硷攻濡炶棄鐣烽锟??�?嬫い鎾跺С缁辨﹢姊绘担鍛婃喐濠殿喚鏁婚獮鎰偅閸愩劎顦梺鍦劋閸ㄧ喖寮告惔銊︾厵闁诡垎鍐╂瘣闂佽�?�掗崢濂革拷?锟介崘顔嘉ч柛鈩兦氶幏褰掓⒑缁嬪潡顎楃痪缁㈠幖椤曘儲绻濋崨顐℃睏闂佸湱鍎ら幐鎾箯缂佹绠鹃弶鍫濆⒔閸掍即鏌熼懞銉х煉鐎殿喗鎮傚畷锟??鍩￠�?顒傛崲閸℃ü绻嗛柣鎰版涧鐢泛鈹戦垾鍐茬殹闁瑰嚖锟???闂佽法鍠曟慨銈咁熆閿燂拷?閺佸啴濡疯缁憋箓鏌ｉ敐鍛伇闁活厽鐟╅幃褰掑箒閹烘垵顬嬪┑鐐靛帶椤﹂潧顫忕紒妯诲�?�缂佸顑欏Λ�?勬⒑缁嬫鍎忔俊顐ｇ箓閻ｇ兘鎮ч崼鐔峰妳闂�?潧绻堥崺鍕洪幖浣瑰仭婵犲﹤鎳庨。濂告偨椤栨侗娈滈柛鈺傜洴楠炴帒螖娴ｅ搫骞堥梺璇茬箳閸嬬喖宕戦幘缁樺剭闁瑰瓨绻嶉悢鍡欐喐鎼达絿鐭欓柟鎹愬煐閿燂拷?????婵＄偑鍊栭崝鎴﹀垂瑜版帪缍栭敓锟???閸曨兘鎷洪柣搴℃贡婵參宕搹鍦＜妞ゆ梻鏅幊鍥煏閸℃洜绐旓�??锟筋噮鍣ｅ畷鐓庘攽鐎ｎ亝鏆梻鍌欒兌缁垶寮婚妸銉殨閻犱浇顫夐敓锟????闂佽法鍠曞Λ鍕Χ缁嬫娼栫紓浣诡焽閿燂�???闂佽法鍣﹂敓�?????????闂佽法鍣﹂敓�?????闂佸憡娲﹂崑鍕磻�?�ュ棛绠鹃悗鐢登瑰瓭濡炪倖鍨甸幊妯虹暦閵夈劊浜归柟鐑樻尵閸樻捇鎮峰⿰鍕煉鐎规洘绮岄埢搴ㄥ箻瀹曞洤骞嬮梻浣侯攰閹活亪姊介崟顖氱９闁绘垼濮ら悡鏇熺箾閸℃绂嬫俊鍙夋尦閺屸槄锟???閿熺瓔鍋嗛幊鍥ㄦ叏婵犲啯銇濓�??锟芥洏鍔嶇换娑㈠箳濠靛懘鍋楁繝纰夋嫹?閿熺晫鍩ｆ鐐寸墵閺佹捇鏁撻敓锟?????婵炶揪绲芥竟濠傤焽閳哄懏鐓犵紒�?�硶娴犳稒绻涢崨顔剧煉婵﹨娅ｉ崠鏍即閻愭祴鎷ら梻浣藉吹閸熸瑩宕堕妸銉ュ⒕闂備礁澹婇崑鍛紦妤ｅ啫缁╅柤鎭掑劘娴滄粓鏌ㄩ悤鍌涘?闂佸搫顑囩划顖滅箔閻斿皝妲堥柕蹇ョ磿閸橀亶鏌熼懝鐗堝涧缂佹煡绠栧鎶筋敆閸曨剛鍘遍梺鍐叉惈椤戝洨寮ч埀顒勬倵鐟欏嫭纾搁柛锟??鍨块妴浣糕枎閹惧磭鐣鹃悷婊冪Ф缁厼顫濋懜纰樻嫽闂佺ǹ鏈悷褔藝閿曞倹鐓欓悹鍥囧懐锛熼梺鐟扮畭閸ㄨ棄鐣烽幒鎴�?敠闁诡垎鍌氼棜婵犳鍠楅敃鈺呭储娴犲纾归柟閭﹀弾濞堜粙鏌ｉ幇顖氱毢缂佺姴顭烽弻鈩冩媴鐟欏嫬纾抽梺璺ㄥ櫐閿燂�??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ょ粣娑㈡煥閻曞倹锟???????闂備線娼чˇ顓㈠磿閺屻儱闂柟鎯板Г閻撴洘銇勯幇闈涗簵闂侇収鍨堕弻锛勪沪閸撗勫垱濡炪�?�鍨哄ú鐔镐繆閸洖宸濇い鏃傛櫕濡差亪姊婚崒娆戭槮缂傚秴锕銊╁�?閻戝棙�?�岄梺鑺ッˇ钘夘焽閺嶃劎绠撅�??锟藉壊鍠曠花浼欐�??閿熻棄鎲＄换鍌炲煘閹达附鍋愰柟缁樺俯娴犲崬鈹戦埄鍐ㄧ祷闁绘鎸搁～蹇撁洪鍕唶闁瑰吋鐣崹濠氬煘濞戞氨纾藉ù锝呮惈鏍￠梺鍦�?濞层倝鎮惧畡鎳婃椽顢旈崟搴涘姂閺佹捇鏁撻敓锟?????缂傚倷绀佹晶搴ㄥ磻閵堝钃熼柣鏂垮悑閻掍粙鏌ㄩ悤鍌涘�??濡ょ姷鍋為敃銏ゅ蓟濞戞ǚ鏋庨煫鍥ㄦ濡箑鈹戦纭锋敾婵＄偠妫勯悾鐑筋敃閿燂拷?�???瀣亜閹烘埊�????閿熶粙宕戦幇顑芥�?闁绘劘灏欓幗鐘电磼椤�?儳校缂佸倸绉撮オ浼村醇椤掍礁�????闂佽法鍠曟慨銈囨崲濠靛鐐婇柤绋跨仛濞呮棃姊婚敓�????閳ь剛鍋涢懟顖涙櫠鐎涙﹩娈介柣鎰絻閺嗘瑩鎽堕弽顓熺厱婵炴垵宕�?▍妯讳繆椤愩垹鏆欓柍瑙勫灴閹瑩寮堕幋鐘辨闂備胶绮�?�鍡椕洪敓锟???閺佹捇鏁撻敓�???????闂備浇顕栭崰妤咃�??锟介崼銉ョ疅闁圭虎鍠栫粈瀣亜閹烘垵浜炴俊鎻掔埣濮婄粯鎷呴崨濠冨枑婵犳鍠氶弫濠氬箖瑜旈幃鈺冩嫚閸欏倶鍎遍湁闁挎繂娲ㄩ妴濠冧繆閹绘帞澧涘ǎ鍥э躬椤㈡盯鎮欙拷?锟芥ɑ娈告俊鐐拷?锟介崑鍕矓閻熼偊娼栨繛宸簻閹硅埖銇勯幘璺轰粶濠碘剝妞藉娲偡閻�?牆鏆堥梺璇�?�枛閸婂潡濡撮敓�????瀵噣宕堕妷銈嗙潖闂備礁�?遍崕銈夊箰閹绢喖绠繛宸簼閳锋垿鏌ｉ幘鍐茬槰婵炶偐鍠栭弻娑欑節閸愨晝顦伴悗娈垮枟閹�?�鐛拷?锟筋喗鍋愰柣銏㈩暜缁卞弶淇婇悙顏庢嫹?閿熻棄顫忔繝姘偍鐟滄棃銆佸Δ鍛潊闁靛牆妫涢崢鎼佹⒑閸涘﹦銆掑褎顨堝☉鍨偅閸愨晜鍤夐梺鍝勭▉閸樹粙鎮￠弴銏＄厵闁煎壊鍓欐俊鑺ョ箾閸涱厽顥炵紒缁樼洴�?�曠厧饪伴崘銊с偖闂佽法鍣﹂敓�?????????闂備胶绮�?�鍥�?磻閿燂拷??闂佸憡鍔︽禍鐐靛婵傚憡鐓犵痪鏉垮船婢ь噣鎮介姘卞煟闁哄苯绉归幐濠冨緞濡儵�?????闂傚倷鑳剁划顖濇懌濡炪�?�姊归悧鐘茬暦閵夆晛宸濋悗娑櫱氶幏缁樼箾鏉堝墽绉繛鍜冪悼閺侇喖鈽夐�?锛勫幈闂�?潧艌閺呮粌鈽夎閹藉爼鎮欙拷?锟藉摜顔曢梺绯曞墲钃遍柟顖氬閺屸剝鎷呴棃鈺勫惈闂佸搫鏈惄顖涗繆閻戣棄绠ｆ繝闈涙处閹烽亶鏌ｆ惔銊︽锭闁活厼鍊搁～蹇撁洪鍜佹濠电偞鍨堕懝楣冿�??锟藉ú顏呪拺缁绢厼鎳忛悵顏堟煕閿燂�??椤ㄥ牓宕氶幒鎾剁瘈婵﹩鍘兼禍閬嶆⒑閸撴彃浜濈紒顔兼捣缁顫濋澶嬪瘜闂侀潧鐗嗗Λ妤佹叏閿曞倹鐓曢悗锝庝簻椤忣參鏌ｅ☉鍗炴珝鐎殿喕绮欓�?�锟??鎮㈢粙鎸庣暯闂傚倷鑳剁划顖炲礉閺囥垺鏅搁柨鐕傛嫹???闂傚倸鍊风粈�???骞栭鈷氭椽濡搁敂钘夊伎闂傚倸鐗婄粙鍫ュ几閿燂拷???/pc闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾婵炶尙鍠栧顐�?磼閻愭潙浠奸柣蹇曞仩濡嫮绮鑸碘拺闁煎鍊曢弸鎴犵磼椤旇偐肖闁告帗甯￠獮妯虹暦閸ャ劍顔曟繝鐢靛Т閿曘�?�宕悩鍙傦綁宕奸妷锔惧帾闂婎偄娲﹀ú鏍ф毄闂備焦鐪归崐鏇灻洪鐑嗘綎婵炲樊浜濋崑锟犳煙濞堝灝鏋欓柧蹇撻叄閺岋絾鎯旈�?鐘叉瘓闂佸憡锕㈢粻鏍春閳ь剚銇勯幒宥堝厡闁哥噦锟?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖宕滆鐢盯鏌涳拷?锟筋煉锟???閿熶粙寮婚敓鐘茬闁靛ě鍐炬毇闂備胶枪鐞氼偊宕濆畝鍕厴闁硅揪绠戠壕鍏肩節婵犲倹�?�呴柟鍑ゆ嫹?闂佽法鍠嶇划娆撳蓟�?�ュ牜妾ㄩ梺鍛婃尪閸斿海鍒掓繝姘鐎规洖娲�?▓楣冩偡濠婂懎顣奸悽顖楁櫊�?�偅绻濋崶銊у帾婵犮垼顕栭崹浼村疮椤栫偞鍊堕柛顐犲劜閳锋垹鐥鐐村櫤闁绘繍浜弻锝呂旈崘銊㈡�?�閻庤娲樺浠嬪极閹剧粯鍋愰柤纰卞墻濡蹭即姊洪懡銈呅ｅù�???绮欏畷婵嬪箣濠㈩亝鐩幃婊堟嚍閵夈垺瀚介梺璺ㄥ櫐閿燂�???????濠电姷鏁搁崑鐐差焽濞嗗緷娲敇閵忊剝娅滈梺缁樺姈濞兼瑧娆㈤悙鐑樼厵闂侇叏绠戞晶浼存煥濞戞艾鏋涙慨濠冩そ楠炲棜顦崇紒鍌氼儔閺屾冻锟???閿熺瓔浜濋崳褰掓煃鐠囪尙效闁诡喒鏅濋幏鐘绘嚑椤掑鏅ｉ梻浣告惈椤︻垶鎮ч崱妯绘珷濞寸姴顑呯粈鍡涙煟閿燂�??閻楀嫭绂嶅⿰鍫熺厪濠㈣埖绋撻悾鍐差熆鐟欏嫸鑰块柡灞界Ф閹叉挳宕熼銈勭礉闁诲氦顫夊ú妯兼暜閹烘缍栨繝闈涱儛閺佸洭鏌ｉ幇顒傛憼闁伙絽銈稿濠氬磼濞嗘帒鍘＄紓渚囧櫘閸ㄥ爼鐛幇顓滃亝闁告劑鍔庨悰銉╂⒑閸濆嫮鈻夐柛妯恒偢閹锋垿鎮㈤崗鑲╁幗闂佸搫鍟导�?�亹閹烘繃鏅梻渚囧墮缁夌敻宕愰崹顐ょ闁瑰鍎愭导鍡涙煙鏉堥箖妾�?柣鎾卞劜閵囧嫰骞樼捄鐑樼亖闂佽法鍣﹂敓锟????闂傚倷绀�?崯鍧楁儍濠靛纾婚柟鍓х帛閸婂爼鏌ｉ幇顒備粵婵炲懏娲栭湁闁绘瑢鍋撻柛銊ョ－濡叉劙骞橈拷?锟芥ê顎撴繛�?�稿Т椤戝懘骞楅悽鍛婄厽闁靛繆鏅涢悘锝夋煕鐎ｎ煉锟???閿熶粙鎮伴敓�????楠炲鏁冮埀顒傜矆鐎ｎ偁浜滈柡宥冨妿閻擃垳绱掗崡鐐靛煟婵﹥妞藉畷銊︾節閸愵煈妲遍梻浣告啞閻熴儵宕幘顔肩畺濞村吋娼欑粻鑽ょ磽娴ｉ�?�姘跺箯缂佹绠鹃柟鐐綑閻掑綊鏌涳�??锟筋偅灏扮紒缁樼⊕閹峰懘宕橀幓鎺戠濠电偛妯婃禍婊冩纯闂備焦鎮堕崕鑽ゅ緤閼恒儳顩查柣鎰靛墯閸欏繑鎱ㄩ敓锟???濡绂嶅⿰鍛亾鐟欏嫭灏俊顐嫹?濠电偛鐗嗛悘婵嗏枍閿燂拷?閺屾冻锟???閿熺瓔浜峰銉╂煥閻曞�?�锟?????婵＄偑鍊戦崹娲偡閳哄懎绠犻柡宥庡幖閻撴稑霉閿濆棗濡抽柡鍥╁亹锟??浠嬫煥濞戞ê顏╁ù婊冦偢閺屾稒绻濋崘顏勨拡闂佽桨绶￠崰妤冩崲濠靛鐐婃い顓熷笚閿燂拷??闂佽法鍠嶇划娆撳蓟閵娾晛鍗抽柣鎴濇处閿燂�???闂佽法鍠撻弲顐ｇ珶閺囥垹閿ゆ俊銈勮兌閸樹粙姊洪崫鍕舵�??閿熸枻锟???閿熺獤鍥х疅闁告縿鍎崇壕濂告煥閻曞倹锟???闂佺ǹ顑嗛幐鎼佸煘閹达附鍋愰柛顭戝亝濮ｅ嫭绻濆▓鍨灍闁圭ǹ鍟块悾鐑藉箛椤斿墽锛滃┑鈽嗗灣缁垶鎮甸悜鑺モ拺闁告繂�?�婵嗏攽閿燂�??椤ユ挻绔熼弴鐔洪檮闁告稑锕﹂崢钘夆攽閻愬弶顥滈柤娲诲灡缁傚秵銈ｉ崘鈹炬嫼闂佺鍋愰崑娑欎繆婵傚憡鐓熼柡宥庡亜鐢埖銇勯弴顏嗙ɑ缂佺粯绻傞～婵嬵敄閳圭偓娅婇柡灞界Ч�?�曨偊宕熼懜闈涱�??闂佽法鍠曟慨銈囩矉�?�ュ鍊烽柣鎴炃氶幏铏圭磽娴ｅ壊鍎愰悗绗涘喛鑰块柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�??????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘绘偘閿燂拷?楠炲鏁冮埀顒傜不濞戙垺鈷掗柛顐ゅ枔閳洘銇勯弬鍨伃婵﹦绮幏鍛村捶椤撶喕寮撮梻浣呵归敃銉╋�??锟芥繝鍌滄殾闁硅揪绠戠粻濠氭偣閸パ冩闁挎洖鍊归悡鏇㈡煛閸ャ儱濡奸柣蹇曞Х缁辨帡鎮╁畷鍥ㄥ垱闂佸搫鏈惄顖烇拷?锟介弴銏℃櫜闁糕剝鐟Σ鐗堜繆閻愵亷锟???閿熻姤顨ラ崫銉х煋闁荤喖鍋婂鏍煣韫囨挻璐￠柣顓熺懄缁绘盯宕卞Ο鍝勫Б闂佸憡鎼╅崜鐔奉潖濞差亜浼犻柛鏇ㄥ墮濞呫�?�绱撴笟鍥ф灍闁瑰摜绮粚杈ㄧ�?閸ャ劌浠虹紓浣割儓濞夋洟藝閺夋娓婚柕鍫濇婢ь剚鎱ㄥΟ绋垮妞ゃ垺鐟︾换婵嬪炊閵娿垺�?�奸梻浣藉吹閸犳劖绔熼崱娑樼闁绘鏁哥壕濂告偣閸ヮ亜鐨洪弽锛勭磽娴ｉ潻�????閿熺晫鏁Δ鍛ч柨婵嗩槸锟??鍐煃閸︻厼浜鹃悗姘偢濮婄粯鎷呯粵瀣秷闂佺ǹ楠搁崥瀣箞閵娾晛围濠㈣泛锕ラ悗顒勬⒒娓氬洤澧紒澶屾暬閹繝寮撮�?锛勫帾婵犵數鍋涢悘婵嬪礉濠婂牊鏅搁柨鐕傛�??????婵＄偑鍊栧褰掝敄濞嗘挸鍚规繛鍡樻尰閻撳啴鏌�?Ο渚▓婵″弶鎮傞幗鍫曟晲婢跺鎷洪梺鍓茬厛閸ｎ噣宕曞☉娆戠闁稿繐鍚嬮埛鎰磼缂佹绠撻柍缁樻崌瀹曞綊顢欓悾灞兼喚濠碉紕鍋戦崐鎴�?礉锟??鍕疇婵せ鍋撴鐐插暢椤﹀磭绱掔紒妯肩疄鐎规洘鍎奸ˇ鎶芥煟鎼搭喖澧ǎ鍥э躬婵℃儼绠涢弴鐐茬厒闂備礁鎽滈崳銉╁垂閸洖绠栭柨鐔哄У閸嬪嫰鏌ゅù�?�珔鐟滄澘瀚板娲箹閻愭彃濮岄梺鍛婃煥缁夎埖绂嶉幖浣哥妞ゆ柨澧介敍婊堟⒑缁嬫寧�?伴柛鎴濈秺�?�曟洟寮�?崼鐔哄幐闁诲繒鍋涙晶浠嬪煡婢舵劖鎳氶柨婵嗩槹閻撴洘绻濋棃娑欘棞妞ゅ繈鍊濋弻鐔虹矙閸喗娈梺璺ㄥ櫐閿燂拷?????闁诲孩顔栭崰鏍偉閻撳海鏆︽繝闈涙閺嬪酣鏌熼幑鎰【缂佷緤绠撻弫鎾绘晸閿燂�??????闂佽法鍣﹂敓�?????????闂備礁鎼ú銊╁磻閻愬樊鍟呮繝闈涱儐閻撶喐绻涢幋婵嗚埞闁哄鐩弻宥囨喆閸曨偆浼岄梺璇″枓閺呯姴鐣疯ぐ鎺濇晝闁挎繂妫涘Σ鎴炵�?閻㈤潧校妞ゆ梹鐗犲畷浼村�?椤撗勬櫔濡炪倖鎸堕崹褰掓倿閸偁浜滈柟鍝勭Ф椤︼箓鏌涢妶搴″⒋闁哄本鐩幃鈺呭箛娴ｅ湱�??????濠电姷鏁搁崑娑樜涘▎鎾崇濠电姵鑹鹃悡鏇㈡煙鏉堥箖妾�?柛�?�剁秮閺屾盯濡烽敐鍛�?�缂備浇灏欑划顖炲Φ閸曨垰绠抽悗锝庝簽娴犻箖姊洪棃娑欐悙閻庢碍婢橀锝夘敋閳ь剟宕洪�?顒併亜閹烘垵顏柛�?�儔閺岋絽螣閸喚姣㈤梺鍝勬４缁犳捇寮婚悢鐓庣濞达絿鍎ら幉锟??姊烘潪鎵槮妞ゆ垵顦靛璇差吋閸偅顎囬梻浣告啞閹稿鎮烽埡鍛畺濡わ絽鍟崐濠氭煢濡警妲烘い鎾存そ濮婅櫣绱掑Ο鍝勵潕闂佽桨鐒﹂幃鍌炲箚閿燂�??瀹曞ジ濡烽敂瑙勫闂備胶顢婇崑鎰板磻濞戙垹绀夋俊銈呮噺閻撴盯鏌涘☉鍗炴灓闁靛棙甯炵槐鎺楊敊绾柉鍚梺杞扮閸熸挳宕洪埀顒併亜閹烘垵顏╅柣鎾达�?�閺�?喐娼忛崜褏鏆犻梺缁樻惈缁绘繈寮诲☉銏犵労闁告劗鍋撻悾鍏肩箾鐎电ǹ袥闁哄懐濮撮～蹇撁洪鍕獩婵犵數濮撮幊搴ㄋ夊┑鍡╂富闁靛牆妫楅悘銉︾箾�?�割喖寮拷?锟芥洩锟???濠碉紕鍋戦崐鏍暜婵犲洦鍤勯柛顐ｆ磸閳ь剨�???????闂備緤锟???閿熻棄鑻晶瀛橆殽閻愬澧柟宄版噹椤垻浠﹂悙�???鏆繝鐢靛Х閺佹悂宕戦悙鍝勫�?�闁诡垱婢樼紞鏃堟⒒娴ｅ憡鎯堟い鎴濇嚇閺屽﹪鏁愭径�?�簵濡炪�?�鍔х粻鎴︽�?�婵犲偆娓婚悗锝庝簼閹癸綁鎷戦柆宥嗏拻濞达絽鎽滈敍宥囩磼椤曞懎鐏︽鐐村姍楠炴牗鎷呴崫銉ュ箣闂備胶顢婇幓顏嗙不閹达附鍋傞柨鐔哄У閻撴洟鏌嶉埡浣告殧濞寸媴濡囩槐鎺楀Ω閵堝洨鐓撳┑顔硷攻濡炶棄鐣烽锟??唯闁靛鍔х紞�???寮婚敐鍛傛梹鎷呴崷顓фЧ闂備焦�?�х换鍕磻閻樼數涓嶆繛鎴欏灩閸楁娊鏌ｅΟ纰辨殰缂佸崬寮剁换婵堝枈濡椿娼戦梺鎼炲妿閺佽鐣烽幋�???绠涢柡澶庢硶閻ゅ洤鈹戦悩缁樻锭妞ゆ垵妫濋崺娑㈠箣閿旇В鎷哄銈嗗姂閸婃洘绂掑⿰鍫熺厾婵炶尪顕ч悘锟犳煛閸涱厾鍩ｆい銏＄懄閹便劑骞囬鍡欐晨濠碉紕鍋戦崐鏍箰妤ｅ啫纾婚柣鎰暩閻岸鏌熺粙璺ㄦ槀濞存粍绮撻弫鎾绘晸閿燂拷???缂傚倸鍊哥粔鎾晝椤忓嫷鍤曞┑鐘崇閸嬪嫮鐥幏�?勫摵闁哄應鏅犲娲濞淬劌缍婂畷鏇㈠蓟閵夈儳顔愰梺褰掑亰閸欏骸鈻撴禒�?�厽闁规澘�???缁ㄥ鏌ｈ箛锝勭盎閼挎劙鏌涢妷鎴濈Х閸氼偊姊虹拠鈥虫灍闁荤啿鏅犻妴�???寮崼婵堫槹濡炪倖鎸荤换鍕涢婊呯＝闁稿本鑹鹃�?顒勵棑缁牊绗熼�?顒勶�??锟介弽顓炲�?�婵炴垶锚閻庮厽绻濋棃娑虫嫹?閿熶粙骞夐敓鐘茬９闁割偅娲橀悡鏇㈡煙娴煎瓨娑ч柡�?�枛閺屽秹鏌�??锟筋亞浼岄梺鍝勬湰缁嬫垿鍩ユ径濠庢建闁割偅绻傞～鐘绘⒒娴ｈ銇熼柛妯煎帶铻炴繝闈涱儏閽冪喖鏌ㄥ┑鍡╂Ц缂佺姵濞婇弻锝夊箛椤旇姤姣勯梺鍝勬閸婃繈骞冮敓�????閳绘捇宕归鐣屼憾闁荤喐绮嶅锟??宕幘顔嘉фい蹇撴噹椤曢亶鏌℃径�?�伌闁哥偛鐖煎铏圭磼濡崵鍙嗛悗娈垮枦椤�?劙骞忛敓�?????闂佽法鍠曞Λ鍕Χ缁嬫娼栫紓浣股戞刊鎾煕濞戞﹫宸ラ柡鍡楃墦濮婃椽鎮烽悧鍫濇殘濠碉�??锟藉级鐢剝淇婇悽绋跨疀闁哄娉曢ˇ銊╂⒑閸愬弶鎯堥柛鐘宠壘鐓ょ紒瀣氨锟??浠嬫煟濡偐甯涙繛鎳峰嫮绠鹃悘鐐诧拷?锟芥俊璺ㄧ磼椤斿墽甯涢柕鍫秮�?�曟﹢鍩￠崘銊ョ疄濠电姷鏁搁崑娑樜涢敓锟???闇夋慨姗嗗墻閻庡墎鎲搁弮鍫濊摕闁靛牆顦痪褔鏌熺粙鍧楋拷?锟藉ù鐘虫尦濮婃椽宕崟顒佹嫳闂佺儵鏅╅崹璺虹暦濞差亝鏅搁柣妯垮皺閿涙粌鈹戦悩璇у伐閻庢凹鍓熷畷瑙勬綇閵娿�?�绠氶梺闈涚墕濞层�?�鏆╅梻浣呵归鍡涙儎椤栫儑�????閿熶粙寮介妸銉х獮闂佸綊鍋婇崜姘舵倵椤掑嫭鈷戠紒�?�硶閻忛亶鏌涳�??锟筋剙鍓抽柟鍑ゆ�??闂佽法鍠撻弲顐ｆ叏閹绢噯�????閿熺晫鎹勯妸�???纾繛鎾村嚬閸ㄨ京鐟ч梻浣筋嚙妤犳悂鎮樺鑸靛亗闁炽儲鍓氬鏍р攽閻樺疇澹樼痪鎯у悑缁绘盯宕卞Ο鍝勵潕闂�?潧鐗婂�???鈥旈崘顔嘉ч柛鈩冾焽椤︺劑姊虹紒姗嗘畼濠殿喗鎸抽幃楣冩倻閽樺娼婇梺闈涚墕濡绂掓總鍛婄厽闊洦娲栨禒褔鏌涳�??锟筋偅灏柍缁樻尰鐎电�?�锟???閿熻姤菤閹锋椽姊洪棃鈺佺槣闁告ê銈稿畷婵撴�??閿熺瓔鍠楅悡娆撴煙闂傚璐版俊顐ｅ灴閺岀喖鐛�?崹顔句紙閻庤娲栧畷顒勶�??锟介崘顏嗙＜婵☆垳绮鎴︽⒒閸屾瑨鍏岄弸顏堟煛閸偄澧伴柛鐘诧工椤撳吋寰勬繝鍕劸闂備胶绮崝妤呭磿閵堝鍋傞柣鏂垮悑閻撴瑩鏌熼鍡楄嫰濞堣泛鈹戦悙鎻掔骇闁瑰憡濞婂濠氭偄绾拌鲸鏅╃紓浣圭☉椤戝棝鎮块敓�????濮婄儤娼幍顔煎闂佸憡姊归悧鐘荤嵁閸℃稑绫嶉柛顐ｇ箘娴煎姊洪懖鈹炬嫛闁告挻鐟╁畷鐢割敆閸曨兘鎷婚梺绋挎湰閻熝囧礉瀹ュ應鏀介柣鎰嚋闊剨�????閿熺瓔鍠撻崝宥咁焽韫囨稑鐓涢柛灞剧⊕椤斿洭姊绘担铏瑰笡闁告梹娲熼幃妯侯潩鐠佸湱绋忛梺鍝勬储閸ㄦ椽鎮�?�▎鎾寸厽闁瑰鍊栭幋鐘辩剨闁规鍠氱壕鏂ゆ�??閿熷鍎遍幊蹇涘窗閿燂拷?閺岋紕浠﹂悙顒傤槰缂備胶绮惄顖氱暦瑜版帩鏁婇柣鎾冲瘨濞笺儵姊绘担钘夊惞濠殿喗娼欑叅闁靛ň鏅涚壕濠氭煏閸繍妲哥紒鐘崇墬娣囧﹪濡堕崨顓熸闂佸摜濮村Λ婵嬪蓟濞戙垹鍗抽柕濞垮劚椤偄顪冮妶蹇氱闁告梹鍨垮濠氭晲婢跺⿴娼婇梺�?�犳〃閼宠埖绂掗銏＄厽闁靛繆鏅涢悘鑼磼缂佹绠烇�??锟筋噮鍋婇獮鍥偋閸績鍋撻柨�?�闁哄鍩堥崕鎰版煥閻曞倹锟???闂傚倷娴囬褔宕欓悾�???�?婇柛鈩冾焽椤╂煡鏌ｉ幇顏囶劅闁轰礁娲弻娑滅�?濮橆兛姹楃紓浣哄█缁犳牕顕ｉ崼鏇為唶婵犻潧妫岄幐鍐磽娴ｅ壊妯堥柛鎾村哺婵＄敻宕熼锝嗘櫇闂�?潧绻嗛弲婊堝煝閸儲鍊垫繛鍫濈仢閺嬫盯鏌涢悢閿嬪仴闁挎繄鍋涜灃闁告侗鍘鹃悿鍕磽娓氬洨鍘滈柟鍑ゆ�??闂佽法鍠撳�???
        .fb_pause({pause_o[2],pause_o[0]}),
        .fb_interrupt(1'b0),       
//        .fb_new_pc(32'b0),
        .new_pc(new_pc_from_ctrl),

        .BPU_flush(BPU_flush),
        .pi_pc1(inst_addr1),
        .pi_pc2(inst_addr2),
        .if_pred_addr1(if_pred_addr1),
        .if_pred_addr2(if_pred_addr2),
        .inst_rreq_to_icache(inst_rreq),
        .pi_is_exception(pi_is_exception),
        .pi_exception_cause(pi_exception_cause),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓顕崑娑⑺夊鑸电厱婵炲棗绻戦幆鍫ユ煃鐟欏嫬鐏撮柟顔规櫊瀹曞綊顢曢敐鍡欐婵犵數濮甸鏍窗濮樿泛绀傛慨妞诲亾濠碘剝鎸冲畷鎺戔槈濮樺吋绁梺璇插嚱缂嶅棙绂嶉悙鏍稿洭顢橀悙鈺傛杸闂佺粯顭囩划顖氣槈瑜庨妵鍕箣濠靛洤娅х紓渚囧枛椤嘲顕ｆ禒�?�垫晣闁绘柨鎼獮鍫ユ⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掞�??锟筋亞鍘介梺闈涳紡閸涱垽绱查梺鑽ゅТ濞层�?�顕ｉ崼�???澶愬閵堝棛鍘搁悗鍏夊亾閻庯綆鍓涜ⅵ婵°�?�濮烽崑娑㈩敄婢舵劕鏋侀柟鐗堟緲瀹告繈鏌涘☉鍗炴灍鐎规洖鐭傞弻鈥崇暆鐎ｎ剛鐦堥悗瑙勬磸閸�?垿銆佸▎鎾崇鐟滃繘宕㈤幒鏃傜＝闁稿本鐟︾粊鏉款渻鐎涙ɑ鍊愭鐐村姈缁绘繂顫濋鍌ゅ數闂備礁鎲＄粙鎴︽偤閵娾晛纾块敓锟???閳ь剛妲愰幒鏂哄亾閿濆簼绨藉ù鐘灮閹叉悂寮堕幐搴闂佸疇顫夐崹鍫曠嵁婵犲洦鐓曞┑鐘插枤濞堟洟鏌熸鏍帨闁瑰嚖锟???闂佽法鍠曞Λ鍕箟閳ュ磭鏆﹂柛娆忣槷缁诲棙銇勯弽銊ф噯妞ゆ帞鍠愮换娑㈠礂閼测晛鈷堢紓浣介哺閹稿骞忛崨�?�樺殐闁斥晛鍟悘锕傛煕閹烘垟搴烽柟鍑ゆ�??闂佽法鍠曞Λ鍕箺濠婂懎顥氶柛蹇氬亹缁犻箖鏌燂�??锟界ǹ鍓冲〒姘洴閺屾稒鎯旈敍鍕唹缂備胶绮惄顖氱暦婵傚壊鏁冮柕蹇曞Х椤旀帞绱撻崒娆愮グ濡炲瓨鎮傞獮鎰節濮橆剛顔嗛梺鍛婄☉閻°劑骞嗛悙鐑樼厽闁绘梻枪椤ュ銇勯幇顑惧仮婵﹦绮幏鍛村川婵犲�?�娈樻繝娈垮枛閿曘�?�绱炴繝鍥ラ柛鎰ㄦ櫇閿燂拷?闂佹悶鍎�?弲娑氱矈閿曞倹鈷戠痪顓炴噺瑜把呯磼閻樺啿鐏撮柨婵堝仱瀹曨煉锟???閿熻姤顭囬崢顏堟⒑閸撴彃浜濈紒璇插暣瀹曠敻宕堕浣哄幈闂佺粯鍔樼亸娆撳春閿濆棙鍙忓┑鐘插暞閵囨繃淇婇銏犳殭闁宠棄顦板蹇涘Ω閹扳晪锟???閿熻棄顫忛搹鍦煓闁割煈鍣崝澶嬬節閻㈤潧浠滈柨鏇樺妼铻為柣鏂款殠濞撳鏌曢崼婵囶棡缁惧墽鏁婚弻娑虫�??閿熺瓔鍋呯亸浼存煙娓氬灝濡界紒缁樼箞瀹曘劑顢氶崨�???鎽嬪┑鐘垫暩閸嬬偤宕硅ぐ鎺戞瀬閻犲洩灏欓弳锕傛煏婵炵偓娅撻柡浣革躬閺屾稖绠涢幘鍗炰划闂佽桨绶℃禍婵堟崲濠靛鍋ㄩ梻鍫熷垁閵夛负浜滈柨婵嗗閻瑩鏌ㄩ悤鍌涘?婵＄偑鍊栫敮鎺楀疮椤栫偞鍋熸い蹇撶墛閻撴瑩鏌涜箛鏇炲付濠殿喖绉归弻鈥崇暆鐎ｎ剛袦闂佽桨鐒﹂崝娆忕暦閸洖惟闁挎梻鏅Σ妤呮⒒閸屾瑦绁版俊妞煎姂閹偤鏁冮崒姘鳖唹闂佹悶鍎洪崜娆撳几閿燂�??閺岀喖宕滆鐢盯鏌￠崨顔斤�??锟介柡宀嬫嫹???闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛鎾茬閸ㄦ繃銇勯弽顐粶缂佺姴缍婇弻宥夊传閸曨剙娅ｇ紒鐐礃椤曆囧煘閹达附鍋愰悹鍥囧嫬�????闂佽法鍠嶇划娆忣嚕閹惰姤鏅濋柛灞剧�?�閸樺崬顪冮妶鍡�?Ё缂佹煡绠栭弫鎾绘晸閿燂拷??闂備浇顕栭崹鎶藉窗閺嶎厼绠栵�??锟藉嫭澹嬮崼顏堟煕閹邦喖浜鹃弫鍫ユ⒒閿燂�??閳ь剚绋撻埞鎺楁煕閿燂�??閸ㄧ敻鎮鹃悜钘夐唶闁哄洢鍔嶉弲銏＄箾鏉堝墽鍒帮拷?锟筋喖澧庨埀顒佷亢閸嬫劗妲愰幘璇茬＜婵炲棙鍩堝Σ顔碱渻閵堝棗鐏ユ俊顐ｇ箞閵嗕線寮�?�閺嬪酣鏌熼幆褏锛嶉柨娑氬枎閳规垿鎮欓弶鎴犱桓闂佸磭顑曢崐婵嬪箖閿燂拷???闂傚倷绀�?幉鈥趁洪敃鍌氬偍濡わ絽鍟崑顏堟煕閺囥劌澧扮紒锟??鍋撶紓浣哄亾濠㈡﹢藝鏉堚晛顥氶柛褎顨嗛悡娑樏归敐鍥╂憘闁搞�?�鐟╅弻锝夋晲閸パ冨箣闂佽鍠撻崹濠氬窗婵犲啯缍囬柕濠忛檮閻濐偄鈹戦悩鎰佸晱闁哥姵顨婇弫鍐煛閸涱厾顦┑鐐叉閹告悂寮搁敓�????閺屾洟宕煎┑鎰ч梺鎶芥敱鐢帡婀�?梺鎸庣箓閹冲繒鎷归敓鐘虫櫢闁跨噦�????婵炲濮撮鍡涙偂閺囥垺鐓忓┑鐐茬仢婵¤姤銇勯妷銉Ч闁靛洤瀚伴、锟??鎮欙�??锟界硶鏁嶉梺璺ㄥ櫐閿燂拷??????闂備礁鎼ú鐘诲礈濠靛鏁傞柣妯款梿瑜版帗鍋戦柛娑卞弾濞差參姊洪悷鏉跨骇闁瑰憡濞婂顐�?箛閺夊灝鑰垮┑鈽嗗灣缁垳娆㈤锔解拻闁稿本鑹鹃�?顒傚厴閹虫宕滄担绋跨亰濡炪倖鐗滈崑娑氱矆婢跺绻嗘い鏍仦閿涚喖鏌ｉ幒鎴敾缂佺粯鐩畷鍗炍熼崫鍕垫綌婵犵數鍋涢幊鎰箾閳ь剚鎱ㄦ繝鍐┿仢妞ゎ澁�????缂傚倷绀�?ˇ閬嶅极婵犳艾绠栭柨鐔哄Т閸楁娊鏌曡箛銉х？闁告﹩浜濈换婵嬫偨闂堟稐绮堕梺璇茬箲缁诲啯绌辨繝鍥ㄥ仼閿燂�??閳ь剙螞椤栨稏浜滈柟鎹愭硾瀛濇繛�?�樼矒缁犳牠寮婚弴銏犵�?�鐟滃秹顢旈鐔翠簻闁靛繆鍓濈粈瀣煥閻曞�?�锟???闂備線娼х换鍫ュ春閸曨垰鑸归柧蹇撴贡绾句粙鏌涚仦鍓ф噭缂佷焦婢橀—鍐级閹寸偞鍠愰梺杞扮贰閸ｏ綁鐛幒锟??鍗抽柣妯跨簿閸╁懘姊婚崒娆愮グ鐎规洖鐏氶幈銊╁级閹炽劍妞芥俊鍫曞川閸屾粌鏋戠紒缁樼箞瀹曟儼顦撮柛鏃撶畱椤啴濡堕崱妤冪憪闂佺粯甯粻鎴︽偩妞嬪簼娌柣鎰靛墮瀵寧绻濋悽闈浶㈤柛鐕佸灦婵￠潧鈹戦幘鏉戭伓?闂佽法鍠曟慨銈吤洪敓�????閵嗗啯绻濋崒銈嗙稁闂佺厧顫曢崐鏇⑺夊鑸碉拷?锟介柨婵嗙凹缁ㄤ粙鏌涢弮鍌涙毈婵﹤顭峰畷鎺戔枎閹烘垵锟???闂備浇顕э�??锟解晝绮欓崼銉ョ柧婵犲﹤鎳忓畷鍙夌箾閹寸偟鎳呯紒�???鍋撻梻浣告啞閸擃剟宕ㄩ婊勬瘞闂傚�?�娴囬褝锟???閿熻В鏅濈划娆撳箳濡炵儵鍋撻敃鍌氱倞闁宠桨�?佽ⅲ闂備緤锟???閿熻棄鑻晶瀛樻叏婵犲啯銇濇鐐寸墵閹瑩骞撻幒鎴綑闂傚�?�绀�?幉锟犲蓟閵娾敡鍥偨閸濄儱绁﹂棅顐㈡处閹峰煤椤忓秵鏅滈梺鍛婁緱娴滄繐锟???閿熻棄銈稿缁樻媴閸涘﹤鏆堢紓浣割儐閸ㄥ潡寮崘顔芥櫆闁告挆鍜冪闯婵犳鍠楁灙闁糕晜鐗犻幃锟犲即閵忕姷顔愬┑鐑囩秵閸撱劑骞忛敓锟????闂佽法鍠嶇划娆忕暦椤愨挌娲敂閸涱垰�?????闂傚倷绀佹惔婊呭緤娴犲缍栭煫鍥ㄦ礈绾惧吋淇婇婵愬殭妞ゅ孩鎹囧娲川婵犲嫧妲堥梺鎸庢磸閸婃繂顕ｉ幎钘夐唶婵犻潧鍟敓�????婵＄偑鍊栧濠氬Υ鐎ｎ亶鍟呴柕澹懐锛濋悗骞垮劚閹锋垿鐓渚囨闁绘劖褰冮弳锝夋煙椤旂晫鐭掗柟绋匡攻缁旂喖鍩為崹顔碱潎闂佸搫鑻粔鐟扮暦椤愶箑绀嬮柤绋跨仛閺嗕即姊绘担鍛婃儓闁瑰嘲顑嗙粋宥夘敂閸曞灚缍庡┑鐐叉▕娴滄粎绮绘导鏉戠閺夊牆澧介幃濂告煟閿濆娑фい顏勫暣婵℃儼绠涢幘鑸敌掗梻浣规偠閸斿宕￠幎鏂ゆ嫹?閿熻棄鈻庨幒鏃傛澑闂佸湱铏庨崹閬嶅棘閳ь剟姊婚敓锟???濞煎骞忛敓�?????闂佽法鍠撻弲顐ょ不閿燂拷???闂傚倸鍊搁崐鐑芥嚄閸撲礁鍨濇い鏍ㄧ箖閹冲矂鏌ｉ悢鍝ョ煁婵犮垺锕㈠畷顖炲箻椤旇�?鍋撻敓锟???瀵噣宕奸锝嗘珖闂備焦瀵у濠氬疾椤愶箑鍌ㄥù鐘差儐閳锋垿鏌熺粙鍨劉缁惧墽鏁婚弻娑虫�??閿熺瓔鍋呭畷�?勬煥閻曞倹锟?????婵犵妲呴崑鍛崲閸繄鏆︽繛宸簼閸婄兘鏌涘┑鍡楊�?妞ゆ挻妞藉娲箰鎼粹懇鎷荤紓渚囧櫘閸ㄨ泛顕ｉ弻銉ョ厸闁告侗鍠掗幏娲煥閻曞倹锟???????闂傚倷鑳舵灙闁挎洏鍎甸獮鎰板箚瑜夐弸搴ㄦ煏韫囧�????閿熶粙宕戦妸鈺傜厱婵炴垶鈽夐崼銉ョ婵炲樊浜濋埛鎴︽煕濞戞﹫鍔熼柍钘夘樀閺屻劑寮村Ο鍝勫Б婵炲瓨绮岄幉鈽呮嫹?閿燂�??锟藉亹閳ь剚绋掗�?�鍥�?储娴犲鈷戦柛鎰�?级閹牓鏌ㄩ弴姗堟嫹?閿熶粙骞冮敓�????閺佸啴宕掑☉姘妇闂備胶纭堕崜婵喢哄⿰鍩跺洭鏁冮崒娑氬帗闁荤姴娲﹂悡锟犲矗閸曨剦娈介柣鎰彧閼板尅锟???閿熻姤娲�?敃銏ゅ箠閻樿鍨傛繛鎴灻兼竟鏇㈡⒑閸撹尙鍘涢柛鐘冲浮瀵劍绂掞拷?锟筋偆鍘介梺褰掑亰閸樼晫绱為幋锔界厽闊洢鍎抽悾鐢告煛锟??瀣М闁诡喓鍨藉鍫曞箣閻樿京�?勫┑掳鍊楁慨鐑藉磻濞戞碍宕叉俊顖濇閺嗭附銇勯幇鍓佺暠閿燂拷?鐎ｎ喗鏅搁柨鐕傛�?????濠电姷顣槐鏇㈠磻閹达箑纾归柡宓本缍庢繝鐢靛У閼瑰墽澹曟繝姘厵闁硅鍔﹂崵娆撴煕濮橆剛绉洪柡灞界Х椤т線鏌涢幘瀵告噰闁糕晝鍋ら獮�?�晜閽樺鍋撻悜鑺ョ厾缁炬澘宕晶顖炴煕閺囥垻鐣烘慨濠呮缁瑩宕犻埄鍐╂毎缂傚�?�娴囬褔鎮ч崱娑欏仼鐎瑰嫭鍣村ú顏嶆晜闁告洦鍘兼慨锔戒繆閻愵亷�????閿熺晫鏁繝鍥ㄢ挃鐎广儱妫涢々鍙夌節婵犲倻澧涢柣鎾寸懇閹鎮介惂鏄忣潐缁傛帡鏁冮崒娑虫�??閿熻姤鎱ㄥ鍡楀箺閿燂拷?鐎ｎ喗鐓涢敓�????閳ь剟宕伴弽褏鏆︽繛鍡樻尭鍥撮梺绯曞墲椤ㄥ繑�?�奸敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏缂佸鍨剁粋鎺撶附閸涘ň鎷哄┑顔炬嚀濞村嫰骞忛敓�?????闂佽法鍠嶇划娆忕暦瑜版帩鏁嗗ù锝勮濞叉悂鎮峰⿰鍛暭閻㈩垱顨婇幃鈥斥枎閹惧鍘介梺鐟邦嚟閸婃牠骞嬮悩杈╁墾闂佹眹鍨归幉锟犳偂閺囥垺鐓涢柛灞剧箖绾爼鏌涢埡�?�М闁哄瞼鍠栭�?�娆戠驳鐎ｎ偆鏆梻浣烘�?瀵爼骞愰幎鑺ユ櫢闁跨噦�??????闂備浇妫勶拷?锟筋剟濡剁粙娆炬綎闁惧繐�?遍惌娆撴煕瑜庨�?�鍛嚕閻楀牏绠鹃悗娑欘焽閻鏌涙惔锝呭付閾荤偤鏌ｉ弬娆炬疇婵炴挸顭烽弻鏇㈠醇濠靛浂妫ゆ繝�???鍥︽喚闁哄本绋撻�?顒婄秵閸嬪棗煤閹绢喗鐓欐い鏇炴閿燂�???闂佽法鍠曡閿燂�??娴犲鍊甸柨婵嗙凹缁ㄨ姤銇勯敓锟???閸旀洟鍩為幋锔斤�??锟介柛銉㈡櫇鏍￠梻浣告啞閹稿鎮烽敂鐣屸攳濠电姴娲﹂崵鍐煃閸濆嫬鏆熼柨娑欑矒濮婅櫣绱掑Ο蹇ｄ邯楠炴牠顢曢敓锟???鐟欙箓鏌涢敂璇插箻缁炬儳銈稿鍫曞醇濞戞ê顬堝┑鐐存儗閸犳濡甸崟顖氼潊闁挎稑瀚崳褔姊猴�??锟界媭鍤欓梺甯秮楠炲啫鈻庨幙鍐╂櫌闂佺ǹ鏈花浠嬪Ψ閳哄�?�鎷绘繛杈剧悼閻℃棃宕靛▎鎾达拷?锟芥繛鎴炲笚濞呭﹪鏌熼搹顐ょ畺闁靛牞缍佸畷锟??濡搁獮顖氭噽绾惧ジ鎮楅敐搴�?�航闁稿簺鍎茬换娑㈠礂閼测晛顫х紓浣虹帛缁嬫垿顢欒箛娑辨晩闁煎鍊曢崵顒勬⒒娴ｈ鍋犻柛濠冪墱閺侇噣鏁撻悩鑼舵憰闂佸搫娲㈤崹褰掓煁閸ャ劎锟??闂傚牊绋掗幖鎰版煛閸涱剛鐭欐慨濠冩そ楠炴劖鎯旈敐鍥╂殼闂備浇顕栭崰鏍ь焽閿熺姴绠栭柣鎴ｆ缁犮儵鏌涢幇顖氱毢濠�?屽灦濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犲ù鐓庣摠閻撴洟鏌熼悜妯诲碍缂佹甯￠弻宥囨嫚閸欏鏀紓浣哄У閻╊垰顕ｉ幘顔藉亜闁告挻褰冮弲顓熺節閻㈤潧啸闁轰焦鎮傞弫鎾绘晸閿燂拷??婵犵數鍋�?崠鐘诲炊閵娿儰缃曢梻浣告啞娓氭宕㈤幖浣歌摕闁挎柨顫曟禍婊堢叓閸ャ劍灏靛褎鐩弻娑虫嫹?閿熺獤鍐ㄢ拤缂備胶绮惄顖氱暦閸楃�?�鐔煎礂閻撳孩鐝紓鍌氾�??锟界粈锟??顢栭崨杈炬嫹?閿熶粙鎮滈挊澶庢憰闂佹寧绻傚Λ娆撳磿閻斿吋鐓忥�??锟界増鐩�?�锕傛惞鎼淬垻锟??婵炲牆鐏濋弸娑㈡煥閺囨ê濡奸柍璇茬Ч閺佹劖寰勬繝鍕瀫闂備礁�?遍搹搴ㄥ窗閺嶎偆鐭嗛悗锝庡亖娴滄粓鏌熸导瀛樻锭濞存粍绻冮妵鍕Ψ閵夘喖鍓伴梺�?�狀潐閸ㄥ潡骞冮埡鍜佹晝闁挎繂鎷嬮埀�???绻樺娲川婵犲啰顦ラ梺璇茬箲锟??鎼佸箖閸ф鏅搁柨鐕傛�??闂佽鍠楅�?�鍛村煝閹捐鍨傛い鏃傛櫕娴滃爼姊绘担铏瑰笡闁圭⒈鍋嗛幑銏犫攽鐎ｎ偄浠掗梺璺ㄥ櫐閿燂�???閻庢鍠曠划娆愪繆閹间焦鏅搁柨鐕傛嫹?濡炪倕�?�╅幑鍥ь潖濞差亝顥堥柍杞拌兌濡诧綁姊洪崨濠庣劷闁告鍥舵晪闁挎繂顦粻锟??鏌ら幁鎺戝姉闁归绮换娑欐綇閸撗呅氬┑鐐叉嫅缁插潡寮灏栨婵炲棙鍨归鏇㈡⒑閸涘﹦鎳冩い锕�?哺閺呭墎鍠婃径�?��??闂佽法鍠曟慨銈吤洪敓�????瀹曟繂顫滈埀顒佷繆閻㈢ǹ绠涢柡澶庢硶椤斿﹪姊虹憴鍕姢闁宦板姂椤㈡棃鎮㈤崗灏栨嫽婵炶揪�???婵倗娑甸崼鏇熺厱闁挎繂绻掗悾鐢告煥閻曞倹锟????????
        .ex_is_bj(ex_is_bj),
        .ex_pc1(ex_pc1),
        .ex_pc2(ex_pc2),
        .ex_valid(ex_valid),
        .real_taken(ex_real_taken),
        .real_addr1(ex_real_addr1),
        .real_addr2(ex_real_addr2),
        .pred_addr1(ex_pred_addr1),
        .pred_addr2(ex_pred_addr2),
        .get_data_req(get_data_req),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠楅悷鈺侇嚕閸洖鍨傛い鏇炴噹濞堫參姊婚崒姘炬�??閿熶粙宕愰幖浣哥９闁绘垼濮ら崐鍧楁煥閺囩儑锟???閿熺晫绮婚弽顓熺厱妞ゆ劧绲鹃敓锟???缂佺偓鍎冲锟犲蓟閿濆绠ｉ柣鎴濇閸斿嘲顪冮妶鍌涙珔鐎殿喖澧庨幑銏犫攽閸モ晝鐦堥梺绋挎湰缁矂路閳ь剟姊绘担鍛佃顨ラ崫銉х煋鐟滅増甯掗拑鐔兼煥濠靛棭妲哥紒鐙呯秮閺岋綁骞囬敓�????閺嗙偟绱掗鑲┬ょ紒顔碱儏椤撳ジ宕ㄩ鍕闂備礁澹婇崑鍡涘窗閹捐鐭楅柛鈩冪⊕閳锋垿鏌涘┑鍡楊仼闁哄棙鐟︾换娑㈠级閹存績鍋撻崹顔炬殾闂傚牊绋堥弸搴ㄦ煙鐎涙ɑ鐓ュù婊呭亾缁绘盯宕煎┑鍫滆檸濠电偛鎳忛敃銏ゅ蓟濞戙垺鏅查煫鍥ㄦ礈琚﹂柣搴㈩問閸犳牠鈥﹂悜钘夊瀭闁诡垎鍛闂佹悶鍎崝宥夋偩閻戣姤鈷戦悹鍥ㄥ絻閸よ京绱撳鍛棦鐎规洘绮岄埥澶娾攦閹冪�?闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊椤掑鏅梺鍝勭▉閸樿偐绮ｅΔ鍛厵闁绘垶锕╁▓鏃堟煟閵堝洤浜剧紒缁樼箖缁绘繈宕掑顓犱壕闂備胶绮敮濠勫垝濞嗘挻鍋傛い鎰剁畱閻愬﹪鏌曟繛鍖℃�??閿熺晫鎹㈤敓�????濮婄儤娼幍顕呮М闂佸摜鍣ラ崹鑸典繆閻㈢ǹ绀嬫い鏍ㄦ皑閿燂拷?闂備礁鐤囧銊╂嚄閼哥數顩峰┑鍌氭啞閳锋帒鈹戦悩鑼闁伙絽鐏氶幈銊︾節閸屻倗鍚嬮悗瑙勬礃鐢帡锝炲┑�?�垫晞闁芥ê顦竟鏇㈡⒑缂佹ê鐏卞┑顔猴�??锟藉畷鐢稿礋椤栨稓鍘遍梺瑙勫礃鐏忔瑩藝閿曞�?�鐓曢柕濠忓缁犳牠鏌曢崶褍顏�??锟筋喕绮欓�?�鏇綖椤撶姵宕熺紓鍌氾�??锟介懗鑸垫叏閹惰棄锟??闁规儼妫勯拑鐔兼煟閺傚灝鎮戦柍閿嬪浮閹鎮介惂鏄忣潐娣囧﹥绂掞�??锟筋�?鎷虹紓浣割儐椤戞瑩宕曡箛鏂讳簻闁瑰瓨绻嶉敓锟???閻庢鍠栭�?�鐑藉箖閵忋倕绀傜痪顓㈡敱閿燂拷??闂佽法鍠曟慨銈夊Φ閸曨垰绠抽柛鈩冦仦婢规洖鈹戦悩顐ｅ�?�閻忕偟鏅禒鎼佹⒑閸濆嫭婀伴柣鈺婂灡娣囧﹪宕奸弴鐐诧拷?锟藉┑鈽嗗灣閳峰牆危瑜版帗鈷掑ù锝呮啞閹牓鏌￠崼顐㈠⒋闁诡垰瀚伴、娑㈡�?�闂堟稓銈﹂梻浣规偠閸庢椽宕滈敃鍌氭瀬闁搞儺鍓氶悡鐔告叏閿燂�??濡寮稿☉妯忓綊鎮崨顖滄殼濠殿喖锕︾划顖炲箯閸涱垳鐭欐繛鍡欏亾椤ユ垿姊绘担鍛靛綊顢栭崱娆愭殰婵°�?�鍟伴惌澶涙�??閿熷鍎遍ˇ浠嬪极閸岀偞鐓曟い鎰剁悼缁犳岸鏌熼懞銉︾闁宠鍨块幃娆撳级閹寸姳鎴烽梻浣虹�?�閺呮冻�????閿熻姤婢�?锝夘敃閿燂�??�???鍐┿亜閺冨�?�娅曢柛姗嗕邯濮婃椽宕滈幓鎺嶇凹缂備浇顕ч崯鏉戠暦閸愯娲敂閸涱垰骞楅梻濠庡亜濞层�?�霉妞嬪海鐜婚柡鍐ｅ亾闁逛究鍔嶇换婵嬪礃閳瑰じ铏庨柣搴ゎ潐濞插繘宕濆鍥ㄥ床婵炴垯鍨圭粻铏�?闂堟稒鍤囬柛瀣殜濮婅櫣鎷犻垾铏亶闂佹寧纰嶉妵鍕敃閿濆洨鐤勫銈冨灪閿曘垽骞冮埡鍜佹晝闁挎繂妫欏▓鐓庘攽閻樺灚鏆╁┑顔惧厴�?�偊宕ㄦ繝鍐ㄥ伎闂佸搫顦伴崵姘洪鍛珖闂佺ǹ鏈銊╂晬濞嗘劒绻嗛柣鎰▕閸庡繒绱掗妸銉у煟鐎规洘鍨块獮妯肩磼濡桨鐢婚梻浣告惈椤︿即顢栧▎寰稑鐣濋崟顑芥嫼闂佸憡绺块崕杈ㄧ墡闂備胶绮〃鍫熸叏閹绢喗鍋╋拷?锟藉嫭澹嬮崼顏堟煕椤愩�?�鏋庡ù婊堜憾濮婃椽宕滈幓鎺嶇凹缂備緡鍠栧ù椋庡垝鐠囧樊娼╅柤鍝ヮ暯閹锋椽姊婚崒姘卞�?缂佸鎸婚弲鍫曞即閻旇櫣顔曢柣蹇曞仜閸嬪﹪骞忛敓�?????闂佽法鍠嶇划娆撳箖瑜庨幆鏃堝Ω閿旇�?�藉┑鐐舵彧缁插潡鎮洪弮鍫濆惞闁告劦鍠楅悡鏇㈡煟濡櫣锛嶅褏鏁搁埀顒冾潐濞叉﹢宕濆▎鎾跺祦闁哄秲鍔嶆刊鎾煟閻旂⒈鏆掗柟顕嗙秮濮婄粯鎷呴搹鐟扮闂佹悶鍔庨崢褑鐏嬮梺鍛婃处閸ㄧ晫绱為弽顓熺厱婵炴垶顭囬幗鐘绘煟閹惧磭绠婚柡灞剧洴椤㈡洟鏁愰崶鈺冩毇闂備線娼婚敓�????濠殿喓鍊濋弫鎾绘晸閿燂拷????闂佹眹鍩勯崹杈╂暜閿熺姴鐏抽柡鍐ㄧ墕�???鍐┿亜閺傛寧顫嶇憸鏃堝蓟濞戙垹鐒洪柛蹇ラ檮锟??鎼佺嵁韫囨梻�???婵﹩鍘搁幏娲⒑閸涘﹦绠撻悗姘煎幗閸掑﹥绺介崨濠勫幈闁诲函缍嗘禍宄邦啅閵夆晜鐓熼柨婵嗘搐閸樻挳鏌ㄩ悤鍌涘?闂備線娼ч悧鍡涘箠鎼达絿鐜绘繛鎴炵懅閿燂拷?闂佹眹鍨藉褍鐡梺璇插閸戝綊宕抽敐澶涙嫹?閿熻棄鈻庨幘鍐插祮闂�?潧楠忕槐鏇㈠储閸涘﹦�???闁靛骏绲剧涵楣冩煥閺囶亪妾柡鍛埣瀵挳鎮滈崱娆忔暩闁荤喐绮岀换妯侯嚕閺屻儺鏁冮柕鍫濇噹閻忓﹪姊洪崫鍕殭闁绘绮撳顐﹀幢濡炴洖缍婇弫鎰板川椤撶噦锟???閿熺晫绱撴担闈涘妞ゆ泦鍥锋�??閿熶粙宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣鍖栭弴鐔哥彅闁诲孩鍑归崜娆忕暤閸曨垱鈷戠憸鐗堝笚閿涚喖鏌ｉ幒鐐电暤闁诡噯绻濋幃銏ゅ礂閼测晛寮虫繝鐢靛█濞佳兾涘▎鎾抽棷閻熸瑥�?�换鍡涙煙缂佹ê淇柣鎾炽偢閺岋�??锟界暆鐎ｎ剛袦闂佽桨鐒﹂崝娆忕暦閸楃偐鏋庨柟瀵稿У濠㈡牠姊虹拠鍙夊攭妞ゎ偄顦叅婵犲﹤鐗嗙粣妤呮煛瀹ュ骸寮块柟鍑ゆ�??闂佽法鍠曞Λ鍕亙闂佸憡渚楅崢楣冩晬濠婂啠�?芥い�???鏋绘笟娑㈡煕閹惧娲存い銏∩戠缓浠嬪川婵炵偓瀚介梺璺ㄥ櫐閿燂�???????闂傚倷鑳剁划顖滄暜椤忓棛涓嶉柟鎯х－閺嗭箓鏌￠崶銉ョ仼閿燂�??閸愵喗鍋″ù锝囨焿閸忓矂鏌熼搹顐ｅ磳闁挎繄鍋涢埞鎴�?醇閻旈锛忛梻浣瑰劤缁绘帒鈻嶉姀銏☆潟妞ゆ洍鍋撴慨濠呮閹风�?骞撻幒鎴炵槪缂傚倸鍊哥粔鏉懳涘┑鍡欐殾闁瑰墎鐡旈敓锟????闁诲孩顔栭崳�???宕戞繝鍌滄殾闁圭儤顨嗛崐鐑芥倵閻㈢櫥褰掔嵁閸喍绻嗛柣鎰典簻閳ь剚鐗犲畷婵嬫晝閸屾氨锛涢梺鍛婃处閸撴艾鈻嶉悩缁樼厵婵炲牆鐏濋弸銈囩棯閹佸仮闁诡喗顨婇弫鎰償濠靛牊鏅肩紓鍌欒兌婵娊宕￠幎钘夎摕鐎广儱娲﹂崰鍡涙煕閺囥劌浜炲ù鐓庣焸濮婅櫣鎷犻垾铏亐闂佸搫鎳忕换鍕ｉ幇鏉跨闁瑰啿纾崰鎰崲濠靛棭娼╂い鎾跺枑椤斿啫鈹戦悩娈挎殰缂佽鲸娲熷畷鎴﹀箣閿燂拷?绾惧綊鏌″搴�?�箹闁搞劌鍊块弻锝夊閳惰泛�?辩划濠氭偐缂佹鍘甸梻渚囧弿缁犳垿宕拷?锟芥ü绻嗛柟缁樺笧婢э箓鏌�?�畝瀣М濠殿喒锟????闂傚倷鑳剁划顖滄暜閹烘鍊舵慨妯挎硾妗呴梺鍛婃处閸ㄦ壆绮婚幎鑺ョ厵閻庢稒顭囩粻銉ッ归悩鑽ょ暫婵﹥妞介獮搴ㄦ嚍閵夛附娈搁梻浣规偠閸斿苯锕㈤崡鐐嶏綁骞囬弶璺啋闁诲孩绋掗敋妞ゅ孩鎸荤换婵嗏枔閸喗鐏嶉梺绯曟櫅閻�?﹦绮嬪鍛�?閻庯綆浜為悿鍕⒑闂堟单鍫ュ疾濞戙垺鍊峰┑鐘插暔娴滄粓鏌熼崫鍕ラ柛蹇撶焸閺屾稑螣閸︻厾鐓撳┑鈽嗗亜閹虫﹢銆�?弴銏�?潊闁炽儲鍓氬Σ閬嶆⒒娴ｅ憡鎯堥悶姘煎亰瀹曟繈骞嬪┑鍫熸濡炪�?�鍔ч梽鍕磹缂佹ü绻嗘い鏍仦濞呮粎绱掗妸銉吋婵﹥妞藉Λ鍐ㄢ槈濮樿京鏆伴梻浣虹�?�閺呮冻�????閿熸垝鍗抽悰顕嗘�??閿熺瓔鍠楅崑鎰版煕閹邦厼绲荤紒銊ｅ劜缁绘繈鎮介棃娑掓瀰濠电偘鍖犻崗鐐洴椤㈡﹢鎮滈崱娆忓Ш闂備礁鍟块幖顐﹀磹閼哥數顩叉繝濠傜墛閻撴瑩鏌熼鍡楄嫰閿燂拷??闂傚倷娴囬褝锟???閿熻В鏅滅粚閬嶅传閸曞孩鐩畷鐔碱敍濮樺崬骞嬮梻浣侯攰閹活亪姊介崟顖氱９闁绘垼濮ら悡鐘绘煙闂傚鍔嶆繛鎳峰嫮绠鹃柟鍐插槻閹虫劗澹曢挊澹濆綊鏁愰崶銊ユ畬缂備浇灏欑划顖滄崲閿燂拷?????闂備椒绱徊鍧楀礂濡警鍤曢柟缁㈠枛椤懘鏌ｅΟ鑽ゅ灩闁告劕澧介崬鐢告煟閻樼儤顏犻悘蹇嬪妼椤斿繘濡烽埡鍌滃幍濡炪�?�鐗楃划灞剧鏉堛劍鍙忓┑鐘插暞閵囨繈鏌＄仦鑺ュ殗闁诡喗鐟╅幊鐘垫崉娓氼垯绱�?繝鐢靛Л閹峰啴宕橀鍛枛闂備緤锟???閿熺晫鈹掗柛鏂跨Ф閹广垹鈹戯拷?锟筋亞顦ㄩ梺宕囨�?閵囨﹢鎼规惔顫箚闁靛牆娲ゅ暩闂佺ǹ顑囬崑銈夊箖瑜旈幃鈺冩嫚閼碱剛鏆繝鐢靛Т閿曘�?�鎮ч崱娑欙拷?锟藉┑鐘叉处閻撳繐鈹戦悙鑼虎闁告梹鎸抽弫鎾绘晸閿燂�?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殘閳ь剙绠嶉崕鍗灻洪妶澶婂瀭婵犻潧娲ㄧ粻楣冩煕閳╁叐鎴犱焊椤撶姷纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍣ｅ畷鐓庘攽閸垺姣囬梻鍌欑閸熷潡骞栭�???鐤い鏍ワ拷?锟介敓锟????闂佽法鍠曟慨銈呯暆閹间礁钃熸繛鎴炃氶弸搴ㄧ叓閸ラ绋诲Δ鏃堟⒒閿燂�??閳ь剛鍋涢懟顖涙櫠婵犳碍鐓曢柟鎹愭硾閺嬪孩銇勯銏㈢閻撱倖銇勮箛鎾村櫣濞寸媭鍙冨娲传閸曞灚笑缂備降鍔戞禍鍫曠嵁閹版澘�?冩い蹇撴閿涙繃绻涢幘纾嬪婵炲眰鍊曢埢宥咁潨閳ь剟寮诲☉銏犖╅柕濠忓閵嗘劕顪冮妶鍡樼┛缂傚秳绀�?锝嗙節濮橆儵銊╂煏婢诡垰鑻弲锝嗙�?閻㈤潧浠╅柟娲讳簽�?�板﹪鎸婃径娑虫�??閿熶粙姊洪敓�????缁夋挳鎯屽Δ鍛厱闁斥晛鍟伴埊鏇㈡煃闁垮鐏╃紒杈ㄦ尰閹峰懘鎯傞崨濠傤�????闂傚倸鍊烽懗鑸电仚闂佹寧娲忛崐鏇㈡晝閵忋倖鐒硷拷?锟姐儱鎳愰崝�???顪冮妶鍡楃瑐闁煎啿鐖煎畷顖炲蓟閵夛妇�??????
        .fb_pred_taken1(fb_pred_taken1),
        .fb_pred_taken2(fb_pred_taken2),
        .fb_pc_out1(fb_pc1),
        .fb_pc_out2(fb_pc2),
        .fb_inst_out1(fb_inst1),
        .fb_inst_out2(fb_inst2),
        .fb_valid(fb_valid),
        .fb_pre_branch_addr1(fb_pre_branch_addr1),
        .fb_pre_branch_addr2(fb_pre_branch_addr2),
        .fb_is_exception1(fb_is_exception1),
        .fb_is_exception2(fb_is_exception2),
        .fb_pc_exception_cause1(fb_pc_exception_cause1),
        .fb_pc_exception_cause2(fb_pc_exception_cause2),
        .fb_instbuffer_exception_cause1(fb_instbuffer_exception_cause1),
        .fb_instbuffer_exception_cause2(fb_instbuffer_exception_cause2)
    );
    wire [1:0] csr_datf;
    wire [1:0] csr_datm;

    wire dcache_is_exception;
    wire [6:0] dcache_exception_cause;

    wire is_tlbsrch;

    reg [31:0] paddr_delayl;
    always @(posedge aclk)
    begin
        if(rst) paddr_delayl <= 32'b0;
        else paddr_delayl <= ret_data_paddr;
    end

    wire [4:0] is_exception_execute1;
    wire uncache_out;

    wire llw_to_dcache;
    wire scw_to_dcache;

    backend u_backend(
        .clk(aclk),
        .rst(rst),

        // from outer
        .is_hwi(intrpt),
        
        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕闈涱潖婵犳艾纾兼繛鍡樺笒閿燂�???闂傚倷鐒︼拷?锟窖兠鸿箛娑樼９婵犻潧顑呴悘鎶芥煥閻曞�?�锟???闂佷紮缍囩换婵嬪蓟閸ヮ剚鏅搁柨鐕傛嫹?濠电偛鐗勯崝鎴濐潖閾忚鍠嗛柛鏇ㄥ亜婵憡绻濆▓鍨灁闁稿﹥绻傞锝夊箵閹哄棗鐗氶梺鍓插亞閸犳捇宕㈡禒�?�拺闁圭ǹ娴风粻鎾绘煙閾忣偄濮嶉柟顔斤�?�閺屽棗顓奸崱娆忓箺??闂備胶绮�?�鍛存晝閿曞倸绠查柕蹇曞Л�???浠嬫倵閿濆骸浜滃ù鐘虫そ濮婂宕掑鍗烆杸闂佽法鍣﹂敓�?????闂備線娼х换鍫ュ磹閺嶎厽鍋傞柡鍥╁亹锟??浠嬫煟濡绲婚柡鍡欏仱閺佹捇鏁撻敓�?????????婵＄偑鍊栧Λ浣规叏閵堝纾归柟閭﹀厴锟??浠嬫⒔閸ヮ剙鏄ラ柡宓苯娈梺璺ㄥ櫐閿燂�????闂佹寧绻傛鍛婃櫠椤旂瓔娈介柣鎰皺婢ф稓绱掔紒妯肩畵闁崇粯鎹囧畷褰掝敊閻ｅ奔鎲鹃梻鍌欑劍鐎笛兠哄澶婄柧闁绘ǹ灏欓弳锔界節婵犲倻澧涢柡鍛箞閺屾稓浠﹂悙顒傛闂佹寧绋撻崰鏍涢崨鎼晝闁靛骏�????閿熺瓔妲遍梻浣告惈閻寰婇崜褏鐭夛�??锟姐儱鎳夐崼顏堟煕閺囨娅冪紒銊ヮ煼濮婃椽宕烽鈩冿�??锟介梺鎼炲妿婢ф寮查崼鏇熷殤妞ゆ帒鍊归敍蹇擃渻閵堝棙灏甸柛�?�枛�?�曟椽鏁愭径瀣幐闂佽法鍣﹂敓锟????闂佸摜濮甸悧鐘荤嵁閸愵喗鍊婚柦妯侯槺妤犲洤鈹戦悙鍙夘棞鐟滄壆鍋ら敓锟???妞ゅ繐妫涚壕浠嬫煕鐏炲墽鎳呴柛鏂跨У閵囧嫰濡搁妷褍鈪甸悗瑙勬磻閸楀啿顕ｉ敓�????????濠电姷鏁搁崑鐐哄垂閸洘鏅濋柍杞扮贰閻掍粙鏌嶉崫鍕舵�??閿熻姤绂嶅⿰鍫熺厵闁告繂瀚ˉ婊兠瑰⿰鍕姢妞ゎ亜鍟存俊鍫曞礃閵娿儱顫撳┑掳鍊楁慨鐢稿箖閸�?偛鏄ラ柣鎰惈缁狅綁鏌ㄩ弮鍥棄濞存粌缍婂娲礈閼碱剙甯ラ梺绋款儏閹冲氦顣鹃梺鍛婃处閸ㄩ亶鍩涢幋鐘电＜閻庯綆鍋掗崕銉╂煕鎼淬垹濮嶉柡宀嬬秮閸┾剝绻濋崒�???妗撻梻浣虹帛娓氭宕板Δ鍐╁床婵犻潧顑呯壕鍏肩�?婵犲倸顏柣锝囧厴濮婄粯鎷呴崨濠傛殘濠电偠顕滅粻鎾崇暦閹达箑�?嬫い鏍ㄧ☉閳ь剙鐏氶妵鍕箻閸楃偟浠鹃梺鎶芥敱閸ㄥ潡寮婚妶澶婄畳闁圭儤鍨垫竟鍕渻閵堝懐绠伴柣鎾愁煼�?�曞爼顢楁担鍝ユ濠电姰鍨奸崺鏍拷?锟介崶锟??�?夐柣鎴ｅГ閳锋垿鏌涘┑鍡楊�?鐞氼亪姊洪崨濠冪叆婵炴挳顥撻崚鎺撶節濮橆剛顦悷婊冾�?瀹曟垿骞樼紒妯轰画闂佸搫顦伴娆徫涘畝鍕拺闁告縿鍎辨牎濠电偛寮剁划鎾诲箠閻愮儤鐒硷�??锟姐儱妫�?▓銉╂⒑闂堟稓澧曢柛濠傛啞缁傚秵銈ｉ崘鈺冨幗闂佺粯鏌ㄩ幖顐︼�??锟芥總鍛婄厱闁绘柨鎼禒褏绱掓潏銊ョ闁归�???閺佹捇鏁撻敓�??????闂佺鍕垫當闁哄嫨鍎甸弻锝夊箛椤掍焦鍎撶紓浣哄�?�缂嶄線寮婚妸鈺佺睄闁搞儺鐓堝Λ鍕箾鐎涙鐭婄紓宥咃工椤繐煤椤忓嫭宓嶅銈嗘尵婵绮敓鐘崇厽闁靛繆鏅涢悘鈩冦亜閵娿儲鍤囬柛鈹垮灲楠炴ê煤缂佹ɑ娅嶉梻浣虹帛椤洭寮幖浣规櫖婵犲﹤瀚换鍡涙煏閸繄绠抽柛鎺嶅嵆閺屾盯鎮ゆ担鍝ヤ桓閻庢鍠栭崯鍧椼偑娴兼潙閱囬柣鏂挎惈楠炴劙姊绘担鍛婂暈濞撴碍顨婂畷鏉款潩椤戠偞妞介獮�???顢欓悾灞藉箞闂備礁鍟块幖顐﹀疮椤愶絿顩烽弶鍫厛濞堜粙鏌ｉ幇顒佲枙闁稿孩妫冮弻鈩冩媴缁嬪簱鍋撻崸�???绠板┑鐘插暙缁剁偤鏌涢埄鍐︿沪濠㈣娲樻穱濠囨�?��?�割喖鍓扮紓浣靛妼閻栫厧鐣烽幋锟??绠荤紓浣姑禒顓㈡⒑閸濆嫷妲规い鎴炵懃铻為敓�????閸曨兘鎷洪梺鍛婄缚閸庤鲸鐗庢俊鐐拷?锟介崝灞轿涘┑鍡╁殨闁哄被鍎卞敮闂侀潧顦崹娲棘閳ь剟姊绘担铏瑰笡闁挎岸鏌ｈ箛鏂垮摵鐎殿喗濞婇崺锟犲川椤�?儳骞堥梺璇插嚱缂嶅棝宕滃▎蹇�?瘎婵犵數鍋涢悺銊у垝鎼淬垻浠氶梻浣哥枃椤曆囨煀閿濆宓佹俊顖濇閺嗭箓鏌涢妷銏℃珔闁绘劕锕濠氬磼濞嗘埈妲梺鍦拡閸嬪棛鍒掗弮鍫濊摕闁靛鍎抽ˇ�???鏌ｆ惔顖滅У闁告挻鑹鹃悾鐑藉蓟閵夛妇鍘遍梺鏂ユ櫅閸熶即鍩婇弴銏＄厽闁规儳顕幊鍛磼鏉堛劍灏伴柟宄版嚇濡啫鈽夊顐ｅ亝闂傚�?�绀�?幖顐︻敄閸℃瑧鐭欓柟鍓х帛閸庡銇勮箛鎾跺缂佺姵姘ㄩ幉闈╂嫹?閿熺瓔鍠栫壕濠氭煏韫囧�????閿熶粙鎮″☉銏℃櫢闁跨噦�????闁诲函缍嗛崜娑溾叺濠德帮�??锟芥慨鐑藉磻濞戞◤娲敇閳ь兘鍋撴担鑲濇棃宕ㄩ鐙呯床婵犵數鍋為崹鍫曟偡閵夆晛鍑犳繛鎴炃氶弨浠嬫煟濡櫣浠涢柡鍡忔櫊閺屾冻�????閿熺瓔鍋嗗ú�?�橆殽閻愯宸ラ柣锝嗙箞瀹曠喖顢曢姀鈶╁亾椤撱垺鈷戦柤鎭掑剭椤忓煻鍥寠婢舵鍔烽梺鍝勭▉閸樹粙鎮￠敐澶屽彄闁搞儯鍔岄崵顒佺箾閸忕厧濮ч柟鍑ゆ�??闂佽法鍠曟慨銈吤洪弽顓勫洭鎮界粙鑳憰闂佸搫娲ㄩ崰鎾剁不妤ｅ啯鐓曟い顓熷灥閺嬫稑鈹戦鑺ョ婵﹨娅ｇ槐鎺懳熼懖鈺冪獥闂備焦鎮堕崝蹇撐涢崟顖ょ稏闊洦鎷嬪ú顏嶆晜闁告侗鍘洪悽濠氭⒒娴ｅ憡鎯堟い锔垮嵆閺佹捇鏁撻敓�???????闂傚倸鍊搁崐鐑芥嚄閸洖绠犻柟鎹愵嚙閸氬綊鏌″搴�?�箹缂佺媴锟?????婵犵數濮烽弫鍛婃叏閻戣棄鏋侀柛娑橈攻閸欏繘鏌熺紒銏犳灍闁稿骸顦…鍧楁嚋闂堟稑顫�?紓浣哄珡閸パ咁啇闁诲孩绋掕摫閻忓浚鍘奸湁婵犲﹤鎳庢禍鎯庨崶褝韬�?┑鈥崇埣瀹曠喖顢�?悙宸拷?锟介梻鍌欑閹诧繝鎮烽妷褎宕叉慨妞诲亾鐎殿喖顭烽弫鎰緞婵犲嫷鍚呴梻浣瑰缁诲�?�螞椤撶倣娑㈠礋椤撶姷锛滈梺璇�?��?�閸愶絾瀵栫紓鍌欑贰閸ｎ噣宕归幎钘夌闁靛繒濮Σ鍫ユ煏韫囨洖啸妞ゆ挻妞藉铏圭磼濡搫顫嶅銈嗘⒐閻楃姴顕ｉ幎鑺ユ櫢闁绘ê鍟块�?顒傛暬閹嘲鈻庤箛鎿冧痪闂佽法鍣﹂敓�?????闂佽�?�╅鏍窗閺嶎厽鍋夊┑鍌氭憸�?�撲線鏌涢鐘插姎閹喖姊洪棃娑辨▓闁哥姵顨堥埀顒勬涧閻�?�寮婚敐澶嬪亹闁告瑥顦遍埞娑㈡�?�濞堝灝鏋熼柟姝屽吹缁晠鎮㈤悡搴�?�祮闂佺粯鏌ㄦ晶搴ｇ不濮樿埖鈷戦梻鍫熺�?�婢ф洘绻涚仦鍌︽�??閿熶粙寮抽埡鍛拻濞达絽鎳欒ぐ鎺濇晞闁糕剝绋掗崕搴€亜閺嶃劍鐨戦柡鍡檮閵囧嫰寮介銏犲闂佽桨�?�?崯鎾蓟閵娾晛妫�?柟绋垮閸庢挻绻涳拷?锟芥鐭婇柛姘儑閹广垹鈽夐�?鐘甸獓闂佺懓鐡ㄧ换鍐磹椤栨埃鏀介柣鎰絻閹垿鏌ｉ悢鍙夋珚鐎殿喛宕甸埀顒婄秵閸犳牠鎮欐繝鍐︿簻闁瑰搫绉烽崗�?勬煕濡湱鐭欐慨濠冩そ�?�曨偊宕熼锝嗩唲闂備胶绮〃鍛存晝椤忓嫷鍤曟い鎰堕檮閻掔�?�锟???閿熷鍎卞Λ娑㈠储娴犲鈷戦梻鍫熺〒婢ф洟鏌熼崘鑼鐎规洜鏁诲畷鍫曞Ω閿燂拷?瀵寧绻濋悽闈浶㈤悗姘煎枤閺侇喖鈽夊杈╋紲濠德帮拷?锟介崯顐�?几閿燂拷???濠碉紕鍋戦崐鏍ь啅婵犳艾纾婚柟鐐暘娴滄粍銇勯幘璺轰沪缂佸本�?�ч妵鍕晝閳ь剛绱炴繝鍥ц摕闁斥晛鍟刊鎾偡濞嗗繐顏╃痪鐐�?▕濮婄儤娼幍顔煎闂佸湱鎳撳ú顓烆嚕椤愶箑绠荤紓浣股戦敓�???????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻娑樷攽閸曨偄濮夐梺绋款儐閹告悂锝炲┑�?�亗閹肩补妲呭楣冩⒒閿燂�??閳ь剛鍋涢懟顖涙櫠椤栫偞鐓熸い鎾楀啯鐝濋悗瑙勬穿缁绘繈鐛惔銊�?癄濠㈠厜鏂傞崕閬嶅Υ閹烘埈娼╅柨婵嗘噸婢规洟鏌ｆ惔銏╁晱闁革綆鍣ｅ畷鎶芥晲閸涱垱娈炬繝闈涳�??锟介幉锟犲磻閸曨垱鐓ｆ慨姗嗗墮閳ь剙顭烽幆鍕償閵婏腹鎷婚梺绋挎湰閻熴劑宕楅敓�?????缂傚倸鍊烽懗鍓佸垝椤栫偛�?夋繛鍡樻尭缁犳岸鏌涢幇闈涙灍闁稿﹤顭烽弻�???螣娓氼垱楔濡炪�?�鏌ㄥΛ娑氭閹捐纾兼繛鍡樺灥婵¤棄顪冮妶搴�?�箹婵炲眰鍔庨崚鎺旂磼濡ǹ浜濋梺鍛婂姂閸斿孩顨ラ崶顒佲拺闁告挻褰冩禍婵堢磼鐠囪�????閿熶粙宕哄☉銏犵睄闁割偆鍠撻崢閬嶆⒑閻熺増鎯堢紒澶嬫綑閻ｇ敻宕卞☉娆戝幐闂佽法鍣﹂敓�?????闂佸摜濮甸幑鍥х暦閻楀牏锟??闁搞儜鍜佹敤闂備胶绮崝鏍ㄧ珶閸℃稑鏋侀柡宥庡幗閳锋帒霉閿濆牆袚闁靛棗鍟扮槐鎺旀媼閸︻厾鐦堥悗瑙勬礃婵炲﹪寮幇鏉垮窛妞ゆ牗绋掗鏇炩攽閻樼粯娑ч柛濠勭帛閻忔瑩姊洪崨濠庢畷濠电偛锕濠氭晲婢跺﹥顥濋梺鍦癸拷?锟解晠宕曢幘婢勬棃鎮╅棃娑楁勃濡炪�?�鍔岄敃銈夛綖韫囨拋娲敂閸曨剙绁舵俊鐐拷?锟介幐楣冨磻濞戞瑤绻嗛柣鎴烆焽閿燂拷?闂佹眹鍨藉褎绂掑⿰鍫熺叆闁哄洦锚閳ь剚绻堥獮鍐箚瑜忛弳瀣煙娴ｅ啯鐝柡鍌�?亾闂傚�?�鑳剁涵鍫曞礈濠靛鍋￠柨鏇�?亾闁崇粯鎹囧鎾閿燂�??閹锋椽姊洪崨濠勨槈闁挎洏鍎甸弫鎾绘晸閿燂�???婵犵數濮幏鍐礃閳哄�?�闂紓鍌欑贰閸犳鎮烽妸褏涓嶆繛鎴欏灩缁犵粯銇勯弽銊�?姇闁哄鎮傚缁樻媴閾忕懓绗″銈庡幖濞层劑宕氶幒妤婃晬婵﹫绲鹃～宥夋偡濠婂啴鍙勫┑锛勬暬瀹曠喖顢涘槌栧悈婵犵數�???濞佳兠洪妶鍛�?�闁靛牆顦伴埛鎴犵磼鐎ｎ亞浠㈤柣锔哄姂閺屾冻�????閿熺瓔浜烽煬顒婃�??閿熺瓔鍠栭�?�鐑藉极閹邦厼绶為悗锝庝簷缁ㄥ姊绘担鍛婂暈缂佸搫娼￠弫鎾绘晸閿燂拷????闂傚倸鍊搁崐鐑芥倿閿燂拷?椤啴宕搁敓�????閸屻劌鈹戦崒婧撳湱澹曡ぐ鎺撶厱鐟滃酣銆冮崼婵堟殼濞撴埃鍋撻柡灞剧洴楠炲洭妫冨☉娆戜憾闂備胶枪閿曪箓宕楅敓�????楠炲啫螖閸涱噮妫冨┑鐐村灦閻燂箓宕伴幇鐗堚拺濞村吋鐟ч悾閬嶆煟濡や焦灏い顐㈢箰鐓ゆい蹇撳椤�?劙姊虹紒妯哄鐟滄澘鍟幈銊ョ暆閸曨兘鎷洪梺鍛婄☉閿曘儵鎮￠妷鈺傗拺閻㈩垼鍠氶崚浼存煟閿濆洤鍘村┑顔瑰亾闂侀潧鐗嗭拷?锟解晠寮插⿰鍫熲拺闁告稑锕ｇ欢閬嶆煕閵婏箑鈻曢柟顖欑窔�?�曞ジ濡烽敂瑙勫婵犳鍠氶幊鎾趁洪妶澶嬶拷?锟介柛娆忣槺缁犳儳霉閿濆懎鏆遍悗姘煎櫍閵嗗懏顦版惔銏犳�?�闂佸搫鍟悧鍡涙嫅閻斿摜绠鹃柟瀵稿仜閻掑綊鏌涳�??锟筋偅宕岄柡浣瑰姈閹棃鍨鹃懠锟??鍤梻浣筋嚙缁绘劕霉濮樿泛鐭楅柛鎰靛枛閽冪噦�????閿熷鍎卞ú锔兼嫹?閿熻姤宀搁弻銈囧枈閸楃偛�???????闂備礁鎼ú锕傛晪婵犳鍠栭崐褰掑Φ閸曨垰顫呴柨娑樺閿燂拷??闂傚倷绀�?幉锛勫垝�???鍕柈闁绘鐗婇崕鐔封攽閻樺弶澶勯柍閿嬪浮閺屾稓浠﹂崜褎鍣梺绋跨箰閻偐妲愰幒妤婃晪闁告侗鍘炬禒鎼佹⒑鐠囷�??锟芥灓闁稿繑锕㈤弫鎾绘晸閿燂�???闂備線娼ч悧鍡涘箠閹扮増鏅繛鎴欏灪閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁梺璇″櫙缁绘繂顕ｉ幘顔碱潊闁挎稑瀚敮鎯р攽閻樺灚鏆╅柛�?�洴閹ê鈹戯拷?锟筋亞顦�?梺闈涚墕椤︿即鎮￠弴銏＄厓闁告繂瀚烽崕鎴︽煙椤旂鍋㈤柡灞界Х椤т線鏌涢幘鏉戝摵妞ゃ垺鐟╁浠嬵敇閻愮儤�?????闁诲氦顫夊ú锟??宕归崜浣瑰床婵犻潧顑呴悙濠囨煃鏉炴媽鍏岄柕鍫檮缁绘繄鍠婂Ο娲绘綉闂佹悶鍔庨弫璇茬暦閹达箑绠涙い鏃傗拡濡粓姊虹粙璺ㄧ婵☆偉娉曢幑銏ゅ幢濡晲绨婚梺鍝勭Р閸斿酣鎯屽畝鍕仺妞ゆ牗绋撻埊鏇㈡煏閸パ冾伂缂佺姵鐩鎾倷鐎甸晲閭┑鐘愁問閸犳牠鏁冮敂鎯у灊妞ゆ牜鍋涚粻顖炴煕濞戞鎽犻柛銈呯Ч閺佹捇鏁撻敓锟????????闂傚倸鍊搁崐椋庢濮橆剦鐒介柤濮愶拷?锟界粈濠囨煕閵夈垺娅囧☉鎾崇Ч閺岀喖骞戦幇闈涙闂佸搫顑勭欢姘跺蓟閻旂厧绀堢憸蹇曟暜濞戙垺鐓涢柛娑卞枟閸婃劙鏌＄仦璇插闁诡噯�?????????
        .new_pc(new_pc_from_ctrl),
        .pc_i1(fb_pc1),
        .pc_i2(fb_pc2),
        .inst_i1(fb_inst1),
        .inst_i2(fb_inst2),
        .valid_i(fb_valid),
        .pre_is_branch_taken_i({fb_pred_taken2,fb_pred_taken1}),
        .pre_branch_addr_i1(fb_pre_branch_addr1),
        .pre_branch_addr_i2(fb_pre_branch_addr2),
        .is_exception1_i(fb_is_exception1),
        .is_exception2_i(fb_is_exception2),
        .pc_exception_cause1_i(fb_pc_exception_cause1),
        .pc_exception_cause2_i(fb_pc_exception_cause2),
        .instbuffer_exception_cause1_i(fb_instbuffer_exception_cause1),
        .instbuffer_exception_cause2_i(fb_instbuffer_exception_cause2),

        .bpu_flush(BPU_flush),   // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷绀�?幉锟犲蓟閵娧呯煋閻犻缚锟??濡插牓鏌ｉ姀鐘冲暈闁稿﹪�?遍妵鍕箣濠靛棛绋忕紓浣靛姀椤曆囷拷?锟介崘顔嘉ч柛鈩冾殔椤洭姊洪幖鐐插鐎规洜鏁搁崚鎺旂磼濡警鍤ら柣搴㈢⊕閿氬ù婊勵殜濮婃椽妫冨☉姘暫濠碘槅鍋勶拷?锟解晝绮嬪鍛牚闁割偁鍨硅ぐ鍕⒑閹肩偛鍔�?柛鏂跨Ф娴滄悂顢橀悢缈犵盎闂婎偄娲ら敃銉モ枍婵犲洦鐓涢敓锟???鐎ｎ剛蓱闂佽鍨卞Λ鍐拷?锟藉▎鎾村亗閹艰揪缍嗛崯鍥�?攽閿涘嫬浜奸柛濞匡拷?锟界粋宥呪堪閸繄鏌堥柣搴㈢⊕鐪夌紒璇叉閺屾盯顢曢敐鍡欘槬濡ょ姷鍋戦崹鐑樼┍婵犲浂鏁嶆繝褏鍋擄�??锟芥稑鈹戦垾铏枙闁告挾鍠庨～蹇曠磼濡顎撻梺缁樺灦閿氭繛鍫濈焸濮婃椽宕妷銉︼拷?锟藉┑鐐碉拷?锟界换婵嗩嚕缂佹锟??闁搞儯鍔嶅▍婊堟⒑閸涘﹣绶遍柛銊ュ船閳绘捇骞嗚�???浠嬫煟濡鍤嬶�??锟芥悶鍎甸弻锝呂旈埀顒勬晝椤忓牆绠栭柣鎰劋閸ゅ啴鏌嶇憴鍕姢濞存粎鍋撻〃銉╂�?�閼碱兛铏庨梺鍛婃⒐绾板秵绌辨繝鍥舵晝闁靛繈鍨婚崝顖毼旈悩闈涗粶缂佺粯鍔楅崣鍛渻閵堝懐绠伴柟鍐差樀楠炲繐煤椤忓應鎷洪梺鍛婄☉閿曪箓鍩ユ径鎰叆闁哄浂浜滈�?�顒傜磼椤旂⒈鐓兼鐐搭焽缁辨帒顫滈崼鐔奉伓?闂佽法鍠曟慨銈夊箞閵娿儙鐔兼偂鎼达拷?锟界帛闁诲孩顔栭崳锟??宕抽敐澶婄濠电姴娲﹂崑鍕煕韫囨艾浜归柛妯圭矙濮婇缚銇愰幒鎴滃枈闂佸摜濮甸〃濠傤嚕閹惰棄鐓涢柛鎰典簼閿涘繘姊虹拠鈥筹拷?锟介柛鎰ㄦ櫅閳ь剦鍨跺娲濞戞瑦鎮欓柣搴㈢濠㈡﹢顢氶敐澶嬫櫢闁跨噦锟???閻庤娲�?崕濂杆囨潏銊�?弿閻熸瑥瀚峰▓婊勬叏婵犲懏顏犵紒杈ㄥ笒铻ｉ柧蹇氼嚃閸庡矂鏌ㄩ悤鍌涘????闁诲孩顔栭崰鏍�??锟介悜钘夋�?�闁圭増婢橀柋鍥煏韫囧鐏繝銏�?�灴濮婄粯鎷呴悜妯烘畬闂佽绻戠换鍫濈暦椤栫儐鏁冮柨鏇楀亾閿燂拷?閸儲鍋ｅΔ锕侊骏閳ь兘鍋撻梺琛″亾闁兼亽鍎禍婊堟煛閸愩劌浜伴柟鍑ゆ嫹?闂佽法鍠嶇划娆忣嚕閵娧呯＜婵☆垰�?辩粻姘舵⒑缂佹ê濮岄柛鈺傜墵钘熷鑸靛姈閻撶喖鏌ㄥ┑鍡樻悙闁告ê鐡ㄩ妵鍕閳╁啰顦伴梺杞扮閸熸挳宕洪�?顒併亜閹烘埊�????閿熶粙鎯岄崱娑欙�??锟介柨婵嗛�?�閺嬬喖鏌ｉ幘�?�樼闁靛洤瀚伴、锟??鎮㈡搴濇樊闂備緤锟???閿熻棄鑻晶鍓х磽瀹ュ嫮绐旓拷?锟筋噮鍋婂畷�???顢欓懖鈺嬬床婵犵數鍋為崹鍓佹暜濡ゅ啠鍋撳顑惧仮婵﹥妞介幊锟犲Χ閸涘懌鍨虹换娑樏癸拷?锟筋偅鐝栨繛瀛樼矌鏋柍璇查叄楠炲鎮╂潏鈺冩喒闂傚倷娴囬崑鎰板煕閸儱�?堟繛鎴炶壘椤ユ艾鈹戦崒姘暈闁稿缍�?弻娑㈠Ψ椤旇崵鐩庨梺姹囧妼閹碱偊鈥﹂懗顖ｆ缂備胶濮甸幑鍥ь嚕婵犳艾鍗抽柕蹇曞Т閼板潡姊洪崫鍕�?窛濠殿喚鍏橀幃浼村閵堝棴锟???閿熻姤绻涢崼婵堜虎婵炲懏锕㈤弻娑㈡晲韫囨洖鍩岄梺浼欑秮锟??杈╃紦娴犲�?堥柛娆忣槹濞呭洭姊绘担鐟邦嚋缂佽鍊歌灋婵炲棙鎸婚崑鐔哥�?闂堟侗鍎愰柍閿嬪浮閺屾稓浠﹂崜褎鍣紓浣瑰姈濮婂湱鎹㈠☉娆愬闁告劖褰冮�?�樼箾閸粎鐭欓柣鎿冨亰瀹曞爼濡搁敂缁㈡О婵＄偑鍊ら崑鍛洪悢鐓庤摕闁跨喓濮撮悙濠囨煏婢跺牆鍔ゅù鐘层偢濮婅櫣绮欓懗顖ｆ蕉闂佸憡姊归崹鍨嚕鐠囨祴妲堟俊顖炴敱椤秴鈹戦绛嬫當闁绘妫欓幈銊モ槈濮樿京锛濇繛杈剧到閹碱偊鍩㈤崼銏㈢＜闁绘ê纾晶顏呫亜閺囶亞绉�??锟芥洖銈稿鎾倷閸濆嫭鏆┑鐘垫暩閿燂�??婵炰匠鍏炬稑鐣濋崟顐ゎ唶闂佸憡鍔︽禍鐐靛閽樺褰掓晲閸涱収妫屽┑鈽嗗灠閻楁捇寮诲☉銏犵闁哄鍨甸幗鍨節绾板纾块柡浣筋嚙閻ｇ兘鎮㈢喊杈ㄦ櫖闂佹寧绻傚Λ娆忊枍閸ヮ剚鈷掑�?�姘ｅ亾婵炰匠鍛床闁糕剝绋戦悿鐐�?婵犲倹鍣介柟鍐叉嚇濮婂宕掑顑藉亾瀹勯偊娓婚柟鐑樻⒐椤洘銇勯敓锟???閸庡磭娆㈤妶鍚ゅ綊鎮╁顔煎壈闁瑰吋娼欓敃顏堝蓟閿涘嫪娌悹鍥ㄥ絻婵洟姊虹粙娆惧剬闁哄懏绮庨幑銏犫攽鐎ｎ偒妫冨┑鐐村灥瀹曨剟宕滄导瀛樷拺缂備焦锚缁楁帡鏌ｈ箛鏂垮摵濠碉紕鏁诲畷鐔碱敍濮�?硸鍞洪梻浣烘�?閻°劎鎹㈠鍡欘浄濠靛倸鎲￠埛鎴犵磽娴ｅ顏嗙箔閹烘鐓熼煫鍥ㄦ煥閸濆搫鈹戦敍鍕毈鐎规洜鍠栭、娑橆潩妲屾牕鏁介梺璇查缁犲秹宕曢崡鐏绘椽鍩￠崘顏嗗箵濠德帮拷?锟介幊蹇涘煕閹达附鐓曟繝闈涘閸�?岸鏌★拷?锟筋亝鎹ｇ紒杈ㄥ笧缁辨帒顫滈崼锝傚亾鐠恒劉鍋撳▓鍨灕妞ゆ泦鍥х叀濠㈣埖鍔曢～鍛存煃閳轰礁鏆為柣婵囧▕濮婅櫣娑甸崨顓濇睏闁荤偞绋忛崕闈涚暦濠婂啠鏀介悗锝庡亜娴犙冣攽閻樼粯娑фい鎴濇�?�曟劙鎮介崨濠備画濠电偛妫楃换鎰邦敂椤忓牊鏅搁柨鐕傛�??闂佸憡鍔︽禍鐐靛閸忕浜滈柡鍐ㄦ搐琚氶悗瑙勬礀閺堫剟銆冮妷鈺傦�??锟介柟缁樺笚閿燂�????闂傚倷绶氬褔鎮ч崱妞㈡稑鐣濋崟顐ゎ唵閻熸粎澧楃敮妤呭煕閹寸姵鍠愰柣锟??鐗嗙粭鎺懨归敓锟???閸楁娊寮诲☉銏�?�亹闁告劖褰冮幗鐢告⒑鐠囷拷?锟芥灓闁稿鎹囨俊鍫曟晲婢跺﹦顦ㄩ梺鍐叉贡閸嬫搫�????閿燂�??锟芥閳规垿鎮欓懜闈涙锭闂佽法鍣﹂敓�??????濠碉紕鍋戦崐鎴﹀磿鏉堚晜宕叉慨妞诲亾鐎殿噯锟??????婵＄偑鍊曠换鎰板箠鎼粹檧鏋嶉柨婵嗩槹閻撶喖鏌熼悙�???鏁鹃柟鍑ゆ嫹?闂佽法鍠嶇划娆忣嚕婵犳艾鐏抽柟棰佺閹垿鏌熼懝鐗堝涧闁瑰嚖�????闂佽法鍠撻弲顐︻敊閿燂拷????闂備浇顫夊畷妯间焊濞嗘垹鐜婚柡鍐ㄧ墛閻撴盯鎮�?悙闈涗壕閿燂�??婢跺瞼纾奸柣妯虹－閳洜绱掔紒妯兼创妤犵偛妫滈ˇ鍗烆熆鐟欏嫭绀嬫慨濠冩そ閹虫牠鍩為悙锟??鐝遍梻浣告啞閹稿鎯勯鐐茬畺闁绘劦鍏欓崑鍛存煕閹般劍鏉归柟椋庣帛缁绘盯骞橀弶鎴犲姲闂佺ǹ顑嗛幐鑽ゆ崲濞戞瑦濯撮柛鎰级婢跺嫰鏌涳�??锟筋亶鍎旈柡灞剧洴閸╁嫰宕橀浣诡潔缂傚倷鑳舵刊顓㈠垂閸洖钃熼柣鏇烇拷?锟介敓锟????闂佽法鍠曟慨銈夛�??锟介崶鈺冧笉闁靛�?濡囩粻楣冩煕韫囨艾浜瑰褜鍓欒彁闁搞儜宥堝惈婵犵锟???閿熺晫鍩ｏ拷?锟芥洏鍔戦�?�锟??鎮㈤崜鎻掓櫃缂傚倸鍊烽懗鍫曞磻閹捐纾块柟鎯版鍥撮梺褰掓？�???�???鎷戦悢鍏肩厽闁哄啫鍊哥敮鍓佺磼閻樺灚鏆柡锟??鍠栭幃婊兾熼懖鈺冩殼闂備礁鎲￠幐缁樼箾婵犲偆娼栭柣鎴灻杈ㄧ箾閸℃ê鐏ラ柛鈺佺焸濮婅櫣鎷犻懠顒傤唹閻庡厜鍋撻柟闂磋兌瀹撲線鏌涢鐘插姎閹喖鏌ㄩ悤鍌涘????闂傚倸鍊烽懗鑸电仚闁荤偞鍑归崑濠傜暦閹邦儵鏃堝川椤撯寬鏇㈡煟鎼搭垳绉甸柛鐘愁殜�?�曟劙鎮介崨濠備画濠电偛妫楃换鎰邦敂椤忓牊鏅搁柨鐕傛�??闂佸憡鍔﹂崰妤呭磻閵婏负浜滈柡宥冨妿閳藉绻涢幖顓炴珝闁哄本鐩崺鐐哄垂椤斿彞鐥梻浣筋嚃閸ㄥ崬螞閸愨晙绻嗛柟闂寸鍞悷婊冪箻瀵爼宕ㄦ繝浣虹畾闂佺粯鍔︽禍鐑藉箯閿燂�???闂佽法鍠嶇划娆忣嚕婵犳艾惟闁宠桨鑳堕鎰渻閵堝棗濮х紒鎻掓健閵嗗懘鎮滈懞銉у幍闂佺粯鍨堕敋闁诲繐绉归弫鎾绘晸閿燂拷??婵炲濮撮鍡涙偂閻旈晲绻嗘い鏍ㄧ箖椤忕姴霉閻樺磭娲撮柡�?嬬節瀹曡精绠涢敓�????閻濇岸鏌ㄩ悤鍌涘�??????婵＄偑鍊栭崝鎴﹀磹閺嶎厼�?嗘繛鎴欏灪閻撱垺淇婇婵嗗惞缂佺姷鍋ら弻锛勪沪缁嬪灝鈷夐悗鍨緲鐎氭悂骞忛敓�?????闂佽法鍠曞Λ鍕櫠鎼达絿鐭氶柛顭戝枓锟??浠嬫煟閹邦剙绾ч柍缁樻�?闇夋繝濠傚缁犵儑锟???閿熻姤娲�?崹鍨暦閻旂⒈鏁冩い鎰剁到閿燂拷????婵＄偑鍊曠换鎰舵�??閿熺晫鍏樺畷婵囧緞婵炵偓�???闂佺粯鍔樼亸娆愭櫠閵忋�?�鐓曢悗锝庡亝鐏忕敻鏌熼獮鍨仼闁宠棄顦甸敓�????闁绘鏁婚悰鎾绘⒒娴ｇ儤�???闁宦板姂閺佹捇鏁撻敓�????????濠电姷鏁告慨鐑藉极閹间礁纾绘繛鎴欏灩鐟欙箓鎮楅敐搴℃灍闁稿绱曢幉姝�?�?濞戞顦梺鍦劋濮婄櫢�????閿熻姤纰嶇换娑㈠级閹搭厼鍓卞銈庡亜缁夌懓顫忓ú顏咁棃婵炴垯鍨诲畷顏嗙磽娴ｄ粙鍝烘繛鑼�?枎閻ｇ兘�???閵堝懎绐涙繝鐢靛Т鐎氼噣鎯�?崼銉︹拺闂傚牊鐩悰婊呯磼閹绘帒鈷旀繛鎴濈仛閵堬綁宕�?埡鍐ㄥ汲闂備礁鎼ù鍌涚椤忓嫷鐎舵い鏂垮⒔绾惧ジ鏌涚仦鍓р槈婵炴惌鍣ｉ弫鎾绘晸閿燂�????闂傚倷绶氬褔鎮ч崱妞㈡稑鈽夐�?鐘插亶闂備緡鍓欑粔鐢稿煕閹达附鈷掗柛顐ゅ枔閵嗘帒顭胯濞叉ɑ绌辨繝鍥舵晝闁挎繂瀛╅悿锟??姊虹拠鈥虫灍闁挎洏鍨藉顐﹀磼閻愯尙顦悷婊冪箻閺佸秴饪伴崨顖滐紳闂佺ǹ鏈悷褔宕濆鍡愪簻妞ゆ挾鍋炲婵堢磼椤旂⒈鐓奸柟顔界懇閹粌螣閻撳骸绠ュ┑锛勫亼閸婃牕螞娴ｅ摜鏆﹂柣銏犳啞閸庢绻涢崱妯哄缂佽妫欓妵鍕箛閳轰胶浠奸梺鍝勬閻熲晛螞娴ｇ懓绶為柟閭﹀幖娴�?垱绻涙潏鍓у埌闁硅绱曢幏褰掓晬閸曨厾锛滄繝銏ｅ煐閿氭繛鍛Ч閺岋拷?锟界暆鐎ｎ剛锛熸繛�?�稿婵″洭骞忛悩瑁佺櫢�????閿熺瓔浜欐竟鏇炩攽閻樼粯娑фい鎴濇噽缁寮介鐔哄幗闂佺鎻徊楣兯夋径�???纾奸柣娆愮懃濞层倗绮昏ぐ鎺擄�??锟芥繛鎴烆伆閹寸姳鐒婂ù鐓庣摠閸婄敻鏌涢�?�鎴濅簽濠⒀嗕含缁辨帗娼忛妸�???纾抽悗瑙勬礃鐢帡鍩㈡惔銊ョ闁挎繂娲ㄥ畷鍫曟⒒閸屾瑧顦﹂柟鑺ョ矋閹便劑鎮介崨濠備罕闂佺粯枪椤曆囨�?�閹惰姤鐓ラ柡鍥╁仜閳ь剙缍婂畷鎰嫚濞村锟??濡炪倖妫佸Λ鍕叏閳ь剟姊虹粙娆惧剱闁圭ǹ顭烽獮蹇涘川椤栨艾顕ч梺鍝勬川閸ｃ儱顭囬弮鍫熲拻濞撴埃鍋撴繛浣冲懏宕查柛鈩冪☉閻掑灚銇勯幒宥囧妽闁诲繘浜堕弻娑虫嫹?閿熺瓔鍋呭畷�?勬煙椤旂晫鐭掗柟绛规�?????闂傚倸鍊烽悞锕傛儑瑜版帒鍨傞悹鍥ㄧゴ閺嬪秹鏌曟径鍫濆Ω濞存粌缍婇弻鐔兼倻濡崵鍙嗙紓浣风筏缁犳垿鍩為幋鐐茬疇闂佺ǹ锕ュú鐔肩嵁婵犲懐锟??婵炴垶顭囬崢閬嶆⒑閸︻厼鍔嬮柛銈嗕亢閵囨劙骞掗幘瀛樼彸闂備礁鎲�?�ú锕傚闯閿燂�??瀹曟繈宕拷?锟芥ǚ鎷洪柣鐐寸▓閳ь剙鍘栨竟鏇炩攽閻愬樊鍤熼柛妯犲洦鍋ら柕濞炬櫆閸嬪�?�绻涢崱妯哄缂佺娀绠栭弻銈嗙附閸撳弶婢撻梺鍝ュ仩濞咃絿妲愰幒锟??惟鐟滃骸鈻嶉弴銏＄厓鐟滄粓宕滃▎鎾达�??锟芥慨姗嗗墻閻斿棝鏌ㄩ悤鍌涘�??闂佽桨绀�?崯鎾拷?锟介弮鍫濈妞ゆ挾鍠愰鏇㈡⒒娴ｇ瓔娼愬鐟版閺呰泛螖閸涱厾锛涢梺绯曞墲椤﹂缚銇愰幒鎾存珳闂佸壊鍋掗崑鍛礊閸儲鈷戝ù鍏肩懆椤撹櫣绱撳鍕槮妞ゎ偄绻戠换婵嗩潩椤掑偊绱叉繝娈垮枟閿曗晠宕楅敓�????瀹曟垿骞樼拠鑼啇婵炶揪绲介幗婊堟晬濞嗘劒绻嗛柣鎰▕閸庡繑绻涳�??锟界ǹ鍘撮柟顖氱焸瀹曞崬螖鐎ｎ偄锟???闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ艾鈹戞幊閸婃鎱ㄩ悜钘夌；闁绘劗鍎ら崑瀣煟濡湱涓查柟鍑ゆ嫹?闂佽法鍠嶇划娆忣嚕閹绢喖顫呴柍鈺佸暞閻濇牠姊婚敓�????閳ь剛鍋涢懟顖涙櫠閹殿喚纾兼い鏃傗拡閻撳ジ鏌熼瑙勬珚闁圭绻濇俊鍫曞川椤撶姴顕遍梻鍌氾拷?锟介悞锕傚箖閸洖纾挎い鏍仜锟??澶愬箹濞ｎ剙濡奸柣鎿勬嫹?閿熺瓔鐔嗛悹楦挎閻忚京鐥幆褋鍋㈤柡宀嬬到铻ｉ柧蹇曟缁辩偞绻濋敓�????閸涱喗姣堥梺鍝勭焿缁辨洘绂掗敃鍌氱鐟滃危閸儲鈷戝ù鍏肩懅缁嬭崵绱掔拠鑼ⅵ鐎规洩�????濠碉紕鍋戦崐鏍暜閹烘柡鍋撳鐓庡濠㈣娲滅槐鎺懳熼懖鈺婂晭闂備胶鎳撻悺銊╂偡閵夆晜鍊舵い蹇撶墛閸婂灚鎱ㄥ鍡�?闁搞�?�娲弻鈥崇暆鐎ｎ剛袦閻庢鍣崜鐔风暦瑜版帩鏁婇柡鍌橈�??锟介敓锟????闂佽法鍠嶇划娆忣潖閾忓湱纾兼俊顖濐嚙閽勫ジ姊虹粙鎸庢崳闁轰浇顕ч锝嗙�?濮橆厽娅滄繝銏ｆ硾閿曘儵藟濠靛鈷戦柛锔诲帎閸︻厸鍋撳☉鎺撴珚鐎规洘娲熼獮妯肩磼濡�?鍋撻崹顐ょ闁瑰鍋熼幊鍛磼閻樻剚鐒界紒杈ㄥ笚濞煎繘濡搁妷锕佺檨闂備浇顕栭崰妤呮偡閳哄拑锟???閿熻棄螖閸涱厾鍔�?銈嗗笒鐎氼剛绮堟径鎰厪闁割偅绻嶅Σ褰掓煟閹惧瓨�?冮柟渚垮妼椤粓宕遍敓锟???閳锋帡姊虹粙鍨劉婵﹤缍婇妴鍐Ψ閳哄偊�????閿熶粙鏌ょ喊鍗炲闁愁亜鐏氱换婵堝枈濡搫鈷夐梺璇�?�枛閸婅绌辨繝鍥ㄧ叆閻庯綆鍋勯崝鍛存⒑闂堟稓绠氭俊鎻掓噹铻為柛鎰靛枟閳锋垹绱掗娑欑闁哄缍婇弻娑虫�??閿熺瓔鍋呯亸顓熴亜椤忓嫬鏆ｅ┑鈥崇埣瀹曞崬螖閸愵亝鍣梻浣筋嚙鐎涒晠宕欒ぐ鎺戠煑闁告劑鍔庨敓�????????婵＄偑鍊曠换瀣倿閿曞�?�鏅搁柨鐕傛�??闂傚倸鍊烽懗鍓佸垝椤栨繃鎳岄柣鐔哥矋濠㈡﹢宕幘顕嗘�??閿熶粙寮�?崼婢冾熆鐠轰警鍎戦柛姗堟嫹???婵＄偑鍊栭崝褏寰婇悾灞芥瀳鐎广儱鎷嬪〒濠氭煏閸繈顎�?ù婊勭箘缁辨帞鎷犻懠锟??鈪靛Δ鐘靛仜閸燁偊鍩㈡惔銊ョ闁告劏鏅滃▍�?勬⒒閿燂�??閳ь剛鍋涢懟顖涙櫠鐎涙ǜ浜滈柕蹇婂墲椤ュ牓鏌ㄩ悤鍌涘�????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠楅悷鈺侇嚕閸洖鍨傛い鏇炴噹濞堫參姊婚崒姘炬�??閿熶粙宕愰幖浣哥９闁绘垼濮ら崐鍧楁煥閺囩儑锟???閿熺晫绮婚弽顓熺厱妞ゆ劧绲鹃敓锟???缂佸墽鍋擄拷?锟窖呮崲濠靛洨锟??闁稿本绮岄�?�娲煥閻曞倹锟???闂佸憡鍔忛弬鍌涚濠婂牏鍙撻柛銉ｅ妽鐏忛潧顭胯濠線骞忛敓�?????闂佽法鍠曟慨銈吤哄Ο鐓庡灊閿燂�??閸曨偆鍘撮梺纭呮彧闂勫嫰寮查鍕厱闁哄洢鍔屾禍妤呮煛婢舵ê寮慨濠呮缁瑩宕犻埄鍐╂毎闂備焦鎮堕崝�?勬�?�濠靛鍋╅柣鎴ｆ閸楁娊鏌曡箛濞惧亾閾忣偒鍚囧┑锛勫亼閸婃牜鏁繝鍕焼濞达綀顫夐崕鐔封攽閻樺弶澶勯柍閿嬪灴閺屾盯骞橀弶鎴犵シ婵炲瓨绮嶇换鍕閹烘梹瀚氶柤纰卞劮閵徛颁簻妞ゆ挾鍋為崰姗堟�??閿熺瓔鍠曠划娆愪繆濮濆矈妲惧銈嗘⒐濞茬喖骞冨Δ鍛仭闁哄顑欏Λ宀勬⒑閸濄儱校婵炲弶绮撻幊鐐烘焼�?�ュ懐顦х紓浣诡殙濡椼劎鑺辨繝姘拺闂傚牊渚楀Σ鍫曟煕鎼淬�?�鐝柡鍛版硾閳藉顫濇潏鈺嬬床缂傚倸鍊烽悞锕傦�??锟介崶顬＄尨�????閿熻姤锕╁▓浠嬫煟閹邦剚鈻曢柛搴㈡閺岀喖顢欓悾灞惧櫘闂佸湱鎳擄�??锟筋厾绮悢纰辨晬婵炴垼椴搁敍鍫濃攽閻樻鏆滅紒杈ㄦ礋�?�曟垿骞嬮敓�????绾惧湱鎲歌箛鎿冨殫濠电姴鍟伴々鐑芥�?�閿濆簼绨芥い锟??鍔曢—鍐Χ閸℃衼缂備胶濮甸崹鍧�?箖閿熺姵鏅搁柨鐕傛嫹?闂佸搫鐬奸崰鎰焽韫囨稑�?堢憸蹇涘汲閻樼粯鈷戠紓浣股戦幆鍫㈢磼缂佹绠烇拷?锟筋喛顕ч埥澶愬閻橀潧濮堕梻浣告啞閸斞呯磽濮橆兘鏌︽い蹇撴绾捐棄霉閿濆娑у┑鈥虫健閺屾稑螣閻樺弶绁柟鍑ゆ�??闂佽法鍠嶇划娆忕暦閿燂拷?椤㈡瑩宕叉竟顖氭处閻撴洟鏌熼幍铏珔濠碉�??锟藉悑閵囧嫰顢楅�?顒勬偋閹炬剚娼栨繛宸簻缁犱即骞栧ǎ锟??鐏╂い锔规櫆缁绘冻锟???閿熻姤顭囬惌銈吤瑰⿰鍕畺缂佸矉�???????婵犵妲呴崹鐢稿磻閹版澘绠犳繝闈涱儐閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曨敊婵劒绨婚梺鍝勬祩娴滅偟绮旈濮愪簻闁靛骏锟???閿熻棄鎽甸梺璺ㄥ櫐閿燂拷??闂佽法鍣﹂敓�??????闂備椒绱徊鍧楀礂閿燂拷?楠炲啴鍩勯崘鈺佸妳濠碘槅鍨崇划顖炲级閹间焦鈷戦悹鍥ㄥ絻閸よ京绱撳鍛棡缂佸倸绉撮埞鎴�??閿熺瓔浜濇潏鍫濐渻閵堝懐绠伴柣锟??锕崺娑㈠箳濡や胶鍘遍柣蹇曞仜婢т粙骞婇崨顔轰簻闁挎棁鍋愰悾鐢告煛閿燂�??閸犳捇宕版繝鍥х闁绘劖澹嗛惄搴ㄦ⒑缂佹ɑ灏柛濠冪箞�?�寮撮悢铏诡啎闂佺粯鍔﹂崜姘舵偟閺冨牊鈷戞慨鐟版搐閳ь兙鍊濆畷鎶芥晲婢跺﹨鎽曞┑鐐村灦缁姴危閻撳寒娓婚柕鍫濆暙婵″ジ鏌熼搹顐㈠闁告帗甯楃换婵嗩潩閸忓吋娅栨繝鐢靛仦閸ㄨ泛顫濋妸鈺婃晩闁哄洢鍨洪崐鐢告煟閻斿憡绶叉い銉ョ箻閺屾盯鎮╅搹顐ゎ槶闂佸ジ缂氭ご鍝ョ紦娴犲宸濆┑鐘插楠炴姊绘担绛嬫綈鐎规洘锚閳绘柨鈽夐�?鐘插殤濠电偞鍨崹娲偂濞戙垺鏅搁柨鐕傛�??闁诲函缍嗛崜娆撳春锟??鍕叄濞村吋鐟х粔�???鏌＄仦鍓р槈闁宠鍨垮畷鍗炍旀繝浣瑰亝缂傚倸鍊烽悞锕傦�??锟�?�箛娑樼煑闁告劦鐓堝鏍ㄧ箾瀹割喕绨奸柛瀣�??锟介獮鏍垝鐟欏嫷娼戝┑鈽嗗亜閺堫剛鎹㈠☉姘ｅ亾濞戞瑯鐒介柣顓滐�??锟介湁婵犲﹤绨肩花缁樸亜閺囶亞鎮奸柟椋庡Т闇夐悗锝庡亽濞兼棃姊婚敓�????濞佳呮崲閹烘挻鍙忛柣銏℃綄婢跺ň鏀介悗锝庡亞閸樹粙姊虹紒妯忣亪宕㈤弽顓熷殝妞ゅ繐鐗婇悡鏇㈡煛閸屾碍鍋ラ柛娆忓閳ь剝顫夊ú妯兼崲閸儻�????閿熻棄鈽夐姀鈽呮�???????婵犵數濮烽弫鎼佸磻濞戙垺鍋嬮柛鈩冪⊕閸婅埖绻濋棃娑卞剰闁告垹�???閺岋綁寮崹顔斤�??锟介梺缁樻尰閻燂箓濡甸崟顖氱睄闁稿本鑹炬禒锟??姊洪柅鐐茶嫰婢ь喗绻涚涵椋庣瘈妤犵偛鍟拷?锟藉ジ骞栭鐔告珦闂傚�?�鐒﹂娆撳垂閻�?牏顩插Δ锝呭暞閻撱儲绻濋棃娑欘棦妞ゅ孩顨婇弻鈽呮嫹?閿熺瓔鍓欓弸娑㈡煛锟??瀣瘈鐎规洏鍔戦、娆撳礈瑜忛崢婊堟⒒娴ｅ憡鎯堥柣顓烆槺缁辩偞绗熼�?�???顕ｉ锟??绠涢柡澶婄仢缁愭盯姊洪崫鍕垫Ч妞ゆ垶鐟︼拷?锟藉ジ宕�?敓锟???缁诲棝鏌曢崼婵囨悙閸熸悂姊虹粙娆惧剳闁稿鍊曢悾宄扳攽閸″繑鐎婚棅顐㈡祫缁插墽绱炴惔銊︹拺闁诡垎鍛啈濡炪�?�鍋勯敓�????闁瑰嚖锟???闂佽法鍠曟慨銈呯暆閹间礁钃熼柣鏃囨绾惧吋淇婇婵囶仩闁荤喆鍔岄埞鎴︻敋閸℃瑧蓱闂佸憡姊归�?�鍫澪ｉ幇鏉跨閻犲洩灏欓敍婊冣攽椤旂即鎴︽儊閻戣棄顫呴柍銉ㄥ皺缁犳艾顪冮妶鍡楀Ё缂佹彃娼￠獮濠囧川椤栨粎锛滃銈嗘⒒閳峰牓宕曡箛鏂讳簻闁规儳鍟块幃鎴嫹?閿熻姤婢橈拷?锟筋厾鎹㈠┑瀣倞鐟滃酣寮抽鍫熲拻闁稿本鐟чˇ锕傛煙绾板崬浜滈悡銈夋煏婵炵偓娅呯紒鎰殜楠炴牕菐閿燂拷?閻忣喗銇勯埡浣哥骇濞ｅ洤锕俊鍫曞川椤斿吋顏￠梻浣瑰▕锟??閬嶅垂閸︻厽顫曢柟铏瑰仦閿燂�???闂佽法鍠撻悺鏃堝储閻ｅ本鍏滈柛鎾茶兌绾惧ジ鏌ｅΟ鍝勬毐闁崇粯娲熼弻锛勪沪閻ｅ睗銏ゆ煟閿濆繒�???妤犵偛绉归�?�娆戝枈鏉堛劍鐦掗梻鍌氾�??锟界粈浣哄椤撶姴鍨濇い鏍仜缁犱即鏌ゆ慨鎰舵嫹?閿熶粙鎯屾径鎰厵闁绘垶蓱閻撴盯鏌涳�??锟筋偅宕岄柡浣瑰姈閹棃鍨鹃懠顒佹櫦闂傚倷绀�?幉锛勬箒缂備緡鍠楅悷銉╋綖韫囨柣鍋婇悷浣碉拷?锟藉Ч妤呮⒑閸︻厼鍔嬮柛銊�?▕�?�曠増绻濋崶銊㈡嫼闂佺鍋愰崑娑欎繆濞差亝鐓曟俊銈勭閳绘洘顨ラ悙鍙夘棦鐎规洘锕㈤�?�娆撴嚍閵夈儱濮冮梻鍌欑窔濞间紮�????閿熻棄鐭傚畷銏°偅閸愨晜娅栧┑鐘诧工閻�?﹪鍩涢幋鐘电＝濞达絽鍘滃Λ銊︺亜韫囨挸鐝嬮柣鏂挎憸閿燂�??闂佹悶鍎崝灞剧濡や胶�???闂傚牊绋戦埀顒佹倐楠炲鏁撻悩鍐蹭簵闂佽法鍣﹂敓�??????闂佺ǹ绻愰ˇ顖涚妤ｅ啯鈷戦梺顐ゅ仜閼活垱鏅讹拷?锟界硶鍋撶憴鍕；闁告鍟块锝嗙鐎ｅ灚鏅ｅ┑鐘欏嫬鍔ゅù婊勫劤闇夐柨婵嗘川閵嗗﹪鏌★拷?锟筋亪鍙勯柡�???鍠栭幃娆擃敆娴ｈ櫣鈻忓┑鐐差嚟婵挳濡堕幖浣哥畺婵°�?�鎳庣粈鍌氼熆鐠虹尨姊楀瑙勬礋濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犻柟缁㈠枟閻撴瑦銇勯弮鍌涘殌濠⒀嗗皺閳ь剙鐏氬姗堟嫹?閿熸垝鍗抽悰�???宕堕澶嬫櫍濠电偞鍨堕悷銉╊敂瑜版帗鈷掗柛灞剧懄缁佸府锟???閿熻姤娲滈弫璇茬暦娴兼潙绠涙い鎾跺Х瑜伴箖姊虹化鏇炲⒉缂佸甯″鏌ヮ敆婵犲啫�????闂佽法鍠庨～鏇㈠磿闁�?单鍥ㄥ鐎涙ê浜楅梺鍝勬储閸ㄦ椽宕愰悽鍛婄叆婵犻潧妫楅弳娆忊攽閳ョ偨鍋㈤柡灞界Х椤т線鏌涢幘鏉戝摵闁诡啫鍏炬棃宕橀鍡欏幇闂佸搫顦悧鍕礉鎼淬劍鏅搁柨鐕傛嫹?闂傚倷鐒﹂幃鍫曞磿椤栫偛�?夐敓�????閸曨偆鍔﹂梺璺ㄥ櫐閿燂拷??濡炪値鍘鹃崗妯侯嚕婵犳艾围濠㈣泛锕﹂悾鎶芥⒑閸︻厼鍔嬮柛銊ョ仛閹便劑寮撮悙鈺傛杸闂佺粯鍔曞鍫曞闯鐟欏嫪绻嗘い鎰剁悼閵嗘帗淇婇崣澶婂妤犵偞顭囬�?顒佺⊕閿氭い搴㈡崌濮婃椽妫冮埡浣烘В闂佸憡顭囨灙閸楅亶鏌涢锝囩婵炴挸顭烽弻鏇㈠醇濠靛浂妫為梺璇茬箞閸庣敻骞冮敓�????椤繈顢曢姀鐘点偖闂佽法鍣﹂敓锟????????婵＄偑鍊栧Λ浣肝涢敓锟????婵犵數濮电喊宥夋偂閻樼粯鐓欐い鎾跺枎缁楁帡鏌涢敓�????椤ㄥ﹪寮婚悢椋庢殝闂侇叏濡囬崥�?�攽椤旂�?�榫氭繛鍜冪悼閸掓帒鈻庨幘宕囶唶闁瑰吋鐣崹鐚存�??閿熻姤濞婂缁樻媴閾忕懓绗�?�┑鈽嗗亜缁绘ê鐣峰⿰鍫熷亜闁兼祴鏅涚粊锕傛椤愩垺澶勭紒瀣浮�?�煡骞栨担鍦�????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺�?喖骞戦幇闈涙闂佹眹鍊楅崑鎾诲Φ閸曨垰绠涢柍鍝勵儐閿燂�???闂佽法鍠嶇划娆忕暦閻熸壋�?介悗锝庡亞閸樺崬顪冮妶鍡�?濠殿喗鎸冲畷婵嗏堪閸喓鍘搁梺鍛婁緱閸犳宕愰幇鐗堢厸閻忕偠顕ф慨鍌炴煙椤旂尨锟???閿熻棄鐣烽幒鎴旀婵妫旈敓锟????婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙盯姊虹紒妯哄闁稿簺鍊濆畷鎴嫹?閿熺瓔鍠楅悡鐔镐繆椤栨繂鍚归敓锟???娴犲鐓冪憸婊堝礂濞戞碍顐芥慨姗嗗墻閸ゆ洟鏌熺紒銏犳灈妞ゎ偄鎳橀弻宥夊煛娴ｅ憡娈插銈呯箳閸犳牕顫忕紒妯诲�?�闁兼亽鍎抽妴濠囨⒑闂堚晝绉剁紒鐘虫崌閺佹捇鏁撻敓锟???????缂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛顐ｆ礀绾惧鏌熼幑鎰靛殭缁炬崘娉曢�?顒冾潐濞叉牕煤閵娧呯焼濠电姴鍊甸弨浠嬫煟濡搫绾ч柟鍏煎姍閺岋箓宕�?鍕拷?锟界紓浣虹帛閻╊垶鐛拷?锟筋亖鏋庨煫鍥ㄦ�?婵爼姊绘担鑺ワ�??锟介敓锟???閿燂�??瀹曨垶骞�?鑹版憰闂侀潧枪閸庮噣寮ㄦ禒瀣厱闁斥晛鍠涙笟娑欎繆椤愮媴锟???閿熶粙鈥旈崘顔嘉ч煫鍥ㄦ皑椤︿即姊虹粙鍧楋�??锟界痪缁㈠幖鍗遍柟鐗堟緲缁犺櫕淇婇妶鍕瓘闁瑰嚖�????闂佽法鍠曟慨銈夊Φ閸曨垰绠抽柛鈩冦仦婢规洟姊绘担鍛婂暈闁哄矉缍佸畷鎰旈崘鈺婃綗闂佸湱鍋撻崜姘跺触鐎ｎ喗鐓曟繝濠傚暙閺嗐垽鏌涘鐓庝喊闁诡喗顨呴埢鎾诲垂椤旂晫浜俊鐐拷?锟介崢楣冨礂濡櫣鏆﹂悷娆忓閸嬪懘鏌涢幇鈺佸闁汇倐鍋撴繝鐢靛仩閹活亞寰婃禒�?�疅闁跨喓濮寸壕瑙勩亜閺嶎偄浠﹂柍閿嬪笒闇夐柨婵嗘噺閸熺偤鏌涢悢鍝勪粶闁靛棙甯掗～婵嬵敇瑜庨悿�???鎮楃憴鍕缂傚秴锕妴浣糕槈濡嘲鐗氶梺鍛婂姂閸斿孩绂嶆导瀛樷拻濞达絽�?卞﹢浠嬫煕閵娿儳绉烘鐐差樀閺佹捇鎮╅崘韫暗闂備胶绮濠氬储瑜忕划鑽ゆ喆閸曨厾顔曢梺鎸庣箓妤犲憡鏅堕敓锟???閺岋�?绠涢敐鍛彎闂佸搫鏈惄顖炲箖閵忋�?�浼犻柕澶堝劚缂佲晠姊绘担鍛婃儓閻炴凹鍋婂畷婵嬪箣閿燂拷?缁犳牠鏌曢崼婵愭Ц缁炬儳鍚嬬换娑㈠箣閻戝洣绶甸梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑缂備胶濮烽崑銈夊箰婵犲洦鍋勯柛蹇氬亹閸橆亪鏌ㄩ悤鍌涘?????闂傚倷鑳剁划顖炲箰婵犳碍鍎庢い鏍仜缁犳牠鏌ㄩ悤鍌涘�??闂佽鍠楅悷鈺呯嵁閹捐绠抽柛鈩兠惁閬嶆⒒閸屾瑧绐�?繛浣冲吘娑樷枎閹寸偞娈伴梺鍦劋椤ㄥ棛绮婚幒妤佲拻濞达綀娅ｇ敮娑㈡煟閻旀潙鍔︽鐐诧躬楠炲洭鎮ч崼婵呮偅闂備焦鐪归崹濠氾拷?锟芥禒�?�；闁规崘鍩栭崰鍡涙煕閺囥劌澧版い锔哄妿缁辨挻绗熼崶褎鐏堢紓浣虹帛鏋俊顐ゅ枎椤啴濡堕崱妯锋嫻闂佹悶鍔嶇换鍕箲閵忋倕骞㈡繛鎴炵懅閸樼數绱撻崒娆戝妽闁挎氨绱掑�???鍠氶悢鍡欐喐鎼粹埗鍝勵潨閳ь剚淇婇悽绋跨妞ゆ牭绲鹃弲婊堟⒑閸涘﹥澶勯柛�?�噹閳绘挾绱掑Ο鑲╃槇闂佽法鍣﹂敓锟?????閻庤娲栧ú銈夋偂閻斿吋鍊甸悷娆忓绾炬悂鏌涢弬鍧�?弰闁糕斁鍋撳銈嗗笒閸婂綊寮抽敓�?????濠电姷顣槐鏇㈠磻濡厧鍨濇繛鍡楁禋濞兼牜绱撴担鑲℃垶鍒婇幘顔界厽闁瑰浼濋鍕ㄦ灁閿燂�??閸曨兘鎷洪梺纭呭亹閸庢垿骞忛敓锟????闂佽法鍠嶇划娆撳箖瑜旈幃鈺呮嚒閵堝懐銈﹂梻濠庡亜濞诧妇绮欓幒�???鐤鹃柟闂寸劍閿燂�????


        .paddr(ret_data_paddr),            // to difftest


        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾婵☆偄鍟悾鐑藉础閻愨晜鐎婚梺瑙勬儗閸ㄨ櫕鎯旀繝鍕＝闁稿本鑹鹃埀顒佹倐�?�曟劙鎮滈懞銉�??閿熶粙鏌ㄩ弴鐐蹭喊闁瑰嚖�????闂佽法鍠嶇划娆忕暦閸洩�????閿熶粙鍩勯崘鈹夸虎濡ょ姷鍋為敃銏わ拷?锟藉▎鎾村仼閻忕偠妫勭粻銉╂⒑鐠囧弶鍞夋い顐㈩槸鐓ら柡宥庣亹濞差亜围濠㈣泛锕﹂崢娲⒑閸撴彃浜為柛鐘叉缁傚秴饪伴崼鐔哄帾闂婎偄娲ら敃銉╋綖婵犲洦鏅搁柨鐕傛�??????闂備礁鎼ú銊╁窗鎼达絿绠旈柟鐑樻尪娴滄粍銇勯幇鍓佹偧缂佺姵鐗楅妵鍕敃閿濆懐浼岄悗娈垮枛閳ь剛鍣ュΣ娲煛婢跺棙娅嗛柨鏇樺灩椤繑绻濆顒傦紲闂佽法鍣﹂敓锟?????闂佸綊妫跨粈浣哄瑜版帗鐓熼柟杈剧到琚氶梺鎼烇拷?锟斤�??锟戒即寮婚妶澶婁紶闁靛闄勫В鍕箾鐎电ǹ校缁炬澘绉电粚杈ㄧ�?閸ヮ煉锟????????闂傚倷鐒﹂幃鍫曞礉鎼淬劌鏋侀悹鍥皺閺嗭附銇勯弽顐粶缂佺嫏鍥ㄧ厵閻庣數枪鏍″┑鐐茬墦缁犳牕顫忓ú顏勪紶闁告洦鍓欓崑宥夋⒑閹肩偛濡芥俊鐐舵閻ｇ兘骞嬮敓锟???鎯熼悷婊冪箻閺佹捇鏁撻敓�????????婵＄偑鍊栭幐楣冨磻濞戞瑦鍙忛柣鎴ｅГ閳锋垹鐥鐐村櫣鐞氭艾鈹戦悙璺虹毢闁哥姴閰ｉ敐鐐剁疀閹句焦妞介�?�鏃堝礋椤撗冩暪闂備胶顢婃竟鍫ュ箵椤忓棗绶ら柛褎顨嗛崑鈺呮⒒閸喍绶辨繛鎾愁煼閺屾洟宕煎┑鍫㈩唶闂佷紮闄勭划鎾诲蓟濞戙垹惟闁靛／鍐幗闂備浇妗ㄩ悞锕傚礉濞嗘挸绠栨繛鍡樻尭娴肩娀鏌涢弴銊ヤ簽闁绘稈鏅犲铏规嫚閹绘帩鍔夌紓浣割儐鐢繝鍨鹃敃鍌氱倞妞ゆ巻鍋撻柛灞诲姂閺岀喖宕滆鐢盯鏌ｉ幘瀵糕槈妞ゎ叀娉曢幑鍕偊閸噮浼冨┑鐐差嚟婵绮婚幋锟??鐓橀柟杈惧瘜閺佸秵绻涢崱妯虹仼闁绘挻鎹囬幃妤冩喆閸曨剛顦ㄥ銈冨妼閻�?﹦绮嬮幒妤佹櫇闁稿本绋戦崜鐟邦渻閵堝棗濮傞柛銊ㄥ吹缁柨煤椤忓懐鍘靛銈嗘⒒閹虫挻鏅堕弻銉︾厵妞ゆ牗绋掗ˉ鍫ユ煥閻曞�?�锟???闂備胶绮敋缁剧虎鍘界粋宥呯暋閹佃櫕�???闂佺粯蓱閸撴岸宕箛娑欑厱闁绘ê纾晶鐢告煛娴ｇǹ鏆ｅ┑锛勫厴婵＄兘顢欓挊澶屾В闂傚�?�娴囨慨銈夋晪濡炪�?�绠撴禍璺侯嚕閹惰姤鏅滃┑顔藉姃缁ㄥ姊虹憴鍕凡濠�?冮叄閹箖鏌嗗鍛板煘濡炪�?�鐗滈崑鐐哄煕閹达附鈷掗柛顐ゅ枍缁惰鲸淇婇幓鎺旂Ш闁哄本鐩顒勬倷閸欏娅ｇ紓浣界堪閸婃洝鐏冮梺鎸庣箓閹冲酣寮冲▎蹇ｆ禆闁告稑鐡ㄩ埛鎴︽煕濞戞﹫�?诲璺哄閺屾盯濡歌椤ｅジ鏌涙惔顔间喊婵﹦绮幏鍛存偡闁箑娈濇繝鐢靛仦瑜板啰绮旈悷鎵殾闁硅揪绠戠粻濠氭煛閸屾ê鍔滈柡鍌�?亾濠碉紕鍋戦崐鏍涢敓锟???瀹曟垿骞囬鐘测叞婵犵绱曢崑鎴�?磹閹达箑�?夊┑鐘叉搐绾惧潡鏌ｉ�?鈶跺湱绮婚弽銊х闁糕剝蓱鐏忎即鏌涢妶鍡楃仸闁靛洤瀚伴獮鎺�?箣濠靛懐鏁栭梻浣告憸閸犲酣顢栨径濠庢綎缂備焦蓱婵挳鏌ら幁鎺戝姷闁瑰嚖锟???闂佽法鍠嶇划娆撳蓟閿濆绠抽柣鎰暩閺嗐倕螖閻橀潧浠﹂柛銊ョ仢閻ｇ兘宕奸弴銊︽櫌?闂備礁鎼鍕濮樿泛钃熼柣鏃傚帶�???鍫㈡喐韫囨洘鏆滄繛鎴欏灪閻撴盯鏌涘☉鍗炴灍闁稿﹥鍔欓弻锛勪沪鐠囨彃顫囬梺璇�?�枔閸婃繂鐣烽幒鎴旀婵妫旈敓锟?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崘鐐暥閻炴碍绻堝缁樻媴閸涘﹤鏆堥梺鍦�?归悥鐓庣暦濠靛绠ｉ柨锟??鍎崇粊锕傛椤愩垺澶勭紒瀣浮�?�煡骞栨担鍦�????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殘閳ь剙绠嶉崕鍗灻洪妶澶婂瀭婵犻潧娲ㄧ粻楣冩煕閳╁喚娈曠紒鍌氼儐缁绘盯宕楅懖鈺侇潷缂備胶绮粙鎴︻敊韫囨侗鏁婇柤濮愶拷?锟介崵顒勬⒒娴ｅ憡鎯堥柟鍐茬箻楠炲啴宕掗悙鑼舵憰闂侀潧艌閺呮粓宕戦崱娑欑厱閻忕偛澧介埥澶愭煥閻曞倹锟????缂傚倸鍊搁崐鎼佸磹閹间礁纾瑰�?�捣閻棝鏌ㄩ悤鍌涘?闁芥ɑ绻冮妵鍕冀椤愩垹澹夐梺杞扮椤戝棝濡甸崟顖氱閻犺櫣娲呴姀銈嗙厱闁靛⿵濡囩粻鎾绘煃鐟欏嫬鐏撮柟顔规櫊�?�曟﹢骞撻幒鎾舵闂傚�?�娴囧銊х矆娴ｈ櫣鐭撶憸鐗堝笒閽冪喖鏌ㄥ┑鍡╂Ц缂佺姵绋掗妵鍕箳閹搭厽笑濠电偛鐗嗛悥鐓庮潖濞差亜宸濆┑鐐搭殘閹虫捁鐏嬮梺鍛婃处閸ㄤ即鎮￠敓锟???閺岀喐娼忛崜褏鏆犻梺缁樻惈缁绘繈寮诲☉銏犵労闁告劗鍋撻悾鍏肩箾鐎电ǹ顎岄柛妯恒偢閳ユ棃宕橀鍢壯囨煕閳╁喚娈樺ù鐘虫倐濮婃椽鎳￠妶鍛瘣闂佸搫鎳忛惄顖炲箖妤ｅ啯鍊婚柤鎭掑労濡啫鈹戦悙鏉戠仸閻㈩垱顨婇幃妤佺節濮橆厸鎷洪梺鑽ゅ枛閸嬪﹪宕甸悢灏佹斀妞ゆ梹鍎抽崢鎾煛娴ｅ摜孝妤楊亙鍗冲畷濂告偄閸欏顏圭紓鍌氾�??锟介崐鐑芥�?�閿曞�?�鏅濋柍鍝勬噺閸婂灝霉閻樺樊鍎愰柣鎾寸☉闇夐柨婵嗘噺閸熺偤鏌熼崣澶嬶�??锟介柡灞稿墲缁楃喖宕惰閻忓牓姊猴拷?锟界姵顥夋い锔炬暬閺佹捇鏁撻敓锟????闂備焦�?�х粙鎴�??閿熺瓔鍓涢弫顔姐偅閸愨斁鎷绘繛杈剧秬椤宕戦悩缁樼厱閹兼番鍨婚惌鎺炴嫹?閿熻姤娲�?敃銏犵暦閿濆唯鐟滃繘鏁嶉悙鐑樷拻濞达絿鐡旈崵娆撴�?�濞戞帗娅婃い銏＄懇瀵粙顢�?悙鐑橈紬??闁诲氦顫夊ú妯荤箾婵犲洤鏋�?柟鐗堟緲瀹告繃銇勯弽銊�?姇妞ゆ梹娲熷缁樻媴缁嬫妫岄梺绋款儏閹冲海鍙呴悗骞垮劚椤︻垶鎮為崹顐犱簻闁瑰搫绉烽崗灞筋熆瑜嶉悘姘跺Φ閸曨垰顫呴柨娑樺閸ｄ即姊洪悷鎵紞闁稿鍊栨穱濠囨�?�閽樺�????????缂傚倸鍊搁崐鎼佸磹閹间礁纾归柣鎴ｅГ閸ゅ嫰鏌涢幘鑼槮闁搞劍绻冮妵鍕�?椤愵�?娌梺绋块�?�鐎涒晠濡甸崟顖氬唨闁靛⿵濡囧▓銈夋⒑閸濆嫭锛旂紒鐘虫崌瀵寮撮悢铏诡啎闂佺粯鍔﹂崜姘舵偟閿曞倹鈷戦弶鐐村椤︼箓鏌涢悢鍛婂唉鐎殿喖顭峰鎾晬閸曨厽婢戦梻浣瑰缁诲倸螞濞戞氨鐜婚柡鍐�??锟界壕钘壝归敐鍕煓闁告繃妞介弻锝夋偆閸屾凹娲梺鐟扮畭閸ㄥ綊鍩為幋�???骞㈤煫鍥ㄦ⒒娴滄牠姊绘担绋款棌闁绘挸鐗撳畷鏉课旈崨顕嗘嫹?閿熶粙鏌涢鐘插姕闁抽攱鍨块弻鐔虹矙閸噮鍔夌紒鍓у亾閹倿寮诲☉娆愬劅闁靛ǹ鍊栭敓�???????闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈咁儐閿燂拷??闂佽法鍠撻弲顐ｆ叏閹绢噯�????閿熺晫鎹勯妸�???纾梺缁樺灦钃遍柟宄板船閳规垿鎮欓懠�???�???闂佺ǹ瀛╂繛濠囧灳閺冨牆绀冩い鏂挎瑜旈弻娑㈠焺閸愮偓鐣堕悶娑滃亹缁辨捇宕掑▎鎺戝帯婵犳鍠氶弫璇茬暦瑜版帒鎹舵い鎾跺仜閻忓﹪姊洪崜鎻掍簮闁瑰啿娲畷鎴﹀箻缂佹ɑ娅滈柟鑲╄ˉ閳ь剝灏欓幐澶娾攽閻愯尙鎽犵紒顔肩Ф閸掓帡骞樼拠鑼舵憰闂佺粯鏌ㄩ崥�?�倿娴犲鏅搁柨鐕傛嫹??闂備礁鎼鍡涙儎椤栫偛钃熼柍钘夋噺閿燂�???闂佽法鍠撻悺�???绂嶉鍫晛婵°�?�鎳忛ˉ鍡楊熆鐠轰警鍎戠紒�???鍋撳┑鐘垫暩婵挳宕愮紒妯绘珷闁靛繈鍊栭悡鐔兼煥濠靛棙顥為柕鍥ㄧ箞閺岋拷?锟界暆鐎ｎ剛锛熸繛�?�稿缁犳挸鐣峰⿰鍡╂Ъ闂佸憡甯楃粙鎴︼拷?锟介崘顔嘉ч柛鎰╁妿娴犳儳鈹戦悙璺虹毢闁哥姵鐗曢锝夘敃閿燂拷?缁犳盯鏌℃径濠勪虎闁兼澘鐏濋埞鎴︽�?�閸欏妫￠柦鍐含閹噣鏁愰崶鈺冿紳闂佺ǹ鏈悢顒勫箯閿燂拷??闂佽法鍠嶇划娆撳箠濡ゅ懎閱囬柡鍥╁仧閿涙盯姊虹憴鍕妞ゆ泦鍛棜闁告牑鍓濋敓锟????闂佽法鍠曟慨銈吤洪弽顬℃椽濡歌閻棗鈹戦悩璇ф嫹?閿熶粙寮ㄦ禒瀣厽婵☆垰鎼痪褔鏌熼崗鐓庡闁哄矉绠撳畷�???顢旈崟顒備邯闂備礁鎼懟顖滅矓瑜版帗鏅搁柨鐕傛嫹???濠电姭鎷冪仦鐣屼桓闂佸搫鏈粙鎴︼綖濠靛鏁嗗璺猴工婢瑰酣姊绘担鍛婃儓闁哄牜鍓涚划娆撳箣閿燂拷?閻擄�??锟筋熆閼搁潧濮囩痪顓涘亾闂備胶绮崝鏇㈠触閳ь剟鏌熼幘顕呮缂佽鲸鎹囧畷鎺戔枎閹达絿鐛ラ梻浣告憸婵�?潧鐣濈粙娆惧殨妞ゆ劧绲块敓锟???濠殿喗锕╅崜婵嬪箺閺囥垺鈷戦柟绋挎捣缁犳挻淇婇锝囨噰鐎规洘娲熼幃銏ゅ礂閼测晛甯鹃梻濠庡亜濞层�?�顢栭崨瀛橈�??锟介柍鍝勬噺閻撴盯鏌涢埥鍡楀箻缂佲檧鍋撴繝娈垮枛閿曘劌鈻嶉敐澶婄闁告洦鍨版儫闂�?潧锟??婵�?�洩銇愬鑸碘拻濞达絿鍎ら敓�????闂佽法鍣﹂敓�?????????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀閹烘娊宕愰弴銏犵柈妞ゆ劧绠戦崹鍌涚節闂堟稒顥戦敓�????娴犲鐓熸俊顖濇閺嬪啫顭跨憴鍕电劷缂佽鲸甯￠幃顏勨枎韫囨梹鎮欑紓浣哄Т缂嶅﹪骞冮敓锟???閳藉鈻嶉搹顐㈢仼濞存粌鎲★�??锟界》锟???閿熻姤顭囬崢鎼佹⒑缁嬫寧�?版い銊ユ噺缁傚秵銈ｉ崘鈹炬嫽闂佺ǹ鏈悢顒勫箯閿燂�???闂佽法鍠嶇划娆撳箠濡ゅ懎�?堝ù锝嚽归悘濠傤渻閵堝棛澧遍柛瀣仱�?�煡顢旈崼鐔哄幗闁瑰吋鐣崺鍕疮韫囨稒鐓曢柣妯虹－婢х敻鏌熼鍝勫姕缂佽桨绮欏畷顐�?Ψ閵壯佸亰闂傚倷绀�?幖顐ょ矙閿燂�??瀹曘垽鎳栭埡鍐х瑝濠电偞鍨崹娲偂閿燂拷???闂備胶绮�?�鍛崲濡櫣鏆﹂柕蹇嬶�??锟介敓锟???闂佺粯鍔忛弲婊堝棘閳ь剟姊洪崷顓炲妺濠电偛锕ら悾鐑藉箛閺夎法顔掗梺鍛婃尫閼冲爼鎮為崗鑲╃闁圭偓娼欓悞褰掓煕鐎ｎ偅宕岄柡灞剧洴閸╃偤宕归鍙ョ礄闁诲孩顔栭崰妤呭箰閹惰姤鏅搁柨鐕傛�??闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡墮閺嬫冻锟???閿熻姤娲�?崹鍧楃嵁閿燂�??瀹曟粍鎷呴搹鐟板Ц婵犵數濮伴崹鐓庘枖濞戙垺鍎旈柤娴嬫櫅椤ユ艾鈹戦崒姘暈闁绘挾鍠愭穱濠囶敍濠靛浂浠╅梺鎸庣☉缁夊綊寮诲澶樻晬婵炴垶鐟чˇ顓犵磽娴ｄ粙鍝洪悽顖滃仧濡叉劙骞掗幊宕囧枛閹虫牠鍩￠崘鈺傜钒闂備浇顕у锕傦綖婢跺⊕鍝勎熼崗鍏兼闂佸湱鍎ら�?�鎰礊閺嶃劎锟??闂傚牊渚楅崕鎰版煛閸涱喚�???闁哄本鐩崺鍕礃閻愵剛鏆柣鐔哥矌婢ф宕曢幎钘夌厴闁硅揪闄勯崑鎰版煕椤垵浜濇慨锝呭缁绘繂鈻撻崹顔界亾闂佺ǹ绻戦敋妞ゆ洩缍�?、鏇㈡晝閳ь剛绮婚悷鎳婂綊鏁愰崨顔藉枑闂佹寧绋掔粙鎴﹀煘閹达附鍊烽柡澶嬪灩娴犙囨⒑閹肩偛濡奸敓�????鏉堚晛鍨濆┑鐘崇閸嬫劗鐥悧鍩亝绂嶆ィ鍐╃厱闊洦鎼╁Σ绋棵瑰⿰鍫㈢暫婵﹥妞藉畷銊︾�?閸愵煈妲遍梻浣呵归鍜冩�??閿熸垝鍗抽獮鍐ㄎ旈崪浣规櫍闂�?潧绻嗗褔骞忓ú顏呪拺闁稿繘妫块懜顏堟煕鎼达紕效妞ゃ垺妫冨畷铏规崉閻戞ê鏋犻梺鍦�?归敃銉ヮ嚗閸曨�?�鐔兼偂鎼粹寬銊╂⒒閸屾瑧顦﹂柟纰卞亞缁瑦绗熼�?�???鐣烽�?锛勵浄閻庯綆鍋勬禍妤呮⒑閹稿海绠撴い锕備憾�?�曪綁骞樼紒妯煎幈闂�?潧锟??缁茶姤淇婃總鍛婄厱闁靛牆楠告晶顖滅磼缂佹娲达拷?锟芥洘顨婇幃鈩冩償閳藉棙缍嶉梻鍌欑窔閳ь剛鍋涢懟顖涙櫠閸欏浜滄い鎰╁焺濡叉悂鎮￠妶澶嬬厸鐎广儱楠哥敮鐐烘煕閵夘喖澧柛�?�ㄥ妿缁辨帪�????閿熺瓔鍘奸崝鐢告煙閼恒儲�?嬫慨濠冩そ�?�曨偊宕熼敓�????缁愭盯姊洪崫銉バｉ柟绋垮⒔閸掓帞绱掑Ο绋夸簼闂佸憡鍔忛弲婵嬪储閸楃儐娓婚柕鍫濋楠炴鏌涢妸褎鏆�??锟筋喚枪閳藉螣闁垮鏉告俊鐐�??锟藉Λ浣规叏閵堝洨鐭嗛悗锝庡亝閸欏繐鈹戦悩鍙夊櫤妞ゅ繒濮风槐鎺撴綇閵娿儳鐟ㄩ柧浼欑秮閺屻�?�霉鐎ｎ偅鐝栫紓浣瑰姈椤ㄥ﹤顫忕紒妯诲�?�閻熸瑥瀚禒鈺呮⒑閸涘﹥鐓ョ紒缁樺姌閻忓姊洪崨濠冨闁搞劎鏅槐鐐哄�?椤撶姴褰勯梺鎼炲劘閸斿酣鍩婇弴銏＄厵妞ゆ牗绮屾禒閬嶆煙椤旂厧妲婚柍璇叉唉缁犳盯骞欓崘褎鍋呯紓鍌欑婢т粙鎼规惔銊ュ瀭閻犺桨�?�?鏍ㄧ箾瀹割喕绨兼い銉ョ墛缁绘稑菐閿燂拷?婵¤偐绱撳鍜冨伐闁伙絿鍏樺鎾閻樼儤鎲伴梻锟??娼ч敓�????缂佺姵鍨剁粋鎺曨樄婵﹥妞藉Λ鍐ㄢ槈濮樿京鏉介梻浣呵归敃銉╂偋閻樿鏄ユ繛鎴欏灩缁狅綁鏌ㄩ弮鍌涙珪闁告ü绮欏铏圭磼濡崵鍙嗛梺纭咁嚋缁辨洖鈻庨�?銈呯煑濠㈣泛鐬奸鏇㈡⒑閸撴彃浜濈痪鏉跨Т閳诲秵绻濋崶銊у幐闁诲繒鍋犻褎鎱ㄩ崒鐐寸厵妞ゆ柨鎼�?顒佺箓閻ｇ兘骞掗幋锟??顫嶅┑顔筋殔濡梻妲愰敓�??????
        .ex_bpu_is_bj(ex_is_bj),
        .ex_pc1(ex_pc1),
        .ex_pc2(ex_pc2),
        .ex_valid(ex_valid),
        .ex_bpu_taken_or_not_actual(ex_real_taken),
        .ex_bpu_branch_actual_addr1(ex_real_addr1),  
        .ex_bpu_branch_actual_addr2(ex_real_addr2),
        .ex_bpu_branch_pred_addr1(ex_pred_addr1),
        .ex_bpu_branch_pred_addr2(ex_pred_addr2),
        .get_data_req_o(get_data_req),
        .csr_dmw0(csr_dmw0),
        .csr_dmw1(csr_dmw1),
        .csr_da(csr_da),
        .csr_pg(csr_pg),
        .csr_plv(csr_plv),

        .asid_in(asid_out),
        .tlbidx_in(tlbidx_out),
        .tlbehi_in(tlbehi_out),
        .tlbelo0_in(tlbelo0_out),
        .tlbelo1_in(tlbelo1_out),
        .tlbehi_out(tlbehi_in),
        .tlbelo0_out(tlbelo0_in),
        .tlbelo1_out(tlbelo1_in),
        .tlbidx_out(tlbidx_in),
        .asid_out(asid_in),
        .ecode_out(ecode_in),
        .rand_index(rand_index),

        .inst_tlb_found(inst_tlb_found),
        .inst_tlb_v(inst_tlb_v),
        .inst_tlb_d(inst_tlb_d),
        .inst_tlb_mat(inst_tlb_mat),
        .inst_tlb_plv(inst_tlb_plv),
        .is_tlbsrch(is_tlbsrch),

        .data_tlb_found(data_tlb_found_out),
        .data_tlb_index(data_tlb_index_out),
        .data_tlb_v(data_tlb_v_out),
        .data_tlb_d(data_tlb_d_out),
        .data_tlb_mat(data_tlb_mat_out),
        .data_tlb_plv(data_tlb_plv_out),
        .invtlb_vpn(invtlb_vpn),
        .invtlb_asid(invtlb_asid),
        .invtlb(invtlb),
        .tlbfill(tlbfill),
        .tlbwr(tlbwr),
        .invtlb_op(invtlb_op),

        .csr_datf(csr_datf),
        .csr_datm(csr_datm),


        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑缂備胶濮烽崑銈夊箰婵犲洦鍋勯柛蹇氬亹閸橆亪鏌ㄩ悤鍌涘?????闂傚倷鑳剁划顖炲箰婵犳碍鍎庢い鏍仜缁犳牠鏌ㄩ悤鍌涘�??闂佽鍠楅悷鈺呯嵁閹捐绠抽柛鈩兠惁閬嶆⒒閸屾瑧绐�?繛浣冲吘娑樷枎閹寸偞娈伴梺鍦劋椤ㄥ棛绮婚幒妤佲拻濞达綀娅ｇ敮娑㈡煟閻旀潙鍔︽鐐诧躬楠炲洭鎮ч崼婵呮偅闂備焦鐪归崹濠氾拷?锟芥禒�?�；闁规崘鍩栭崰鍡涙煕閺囥劌澧版い锔哄妿缁辨挻绗熼崶褎鐏堢紓浣虹帛鏋俊顐ゅ枎椤啴濡堕崱妯锋嫻闂佹悶鍔嶇换鍕箲閵忋倕骞㈡繛鎴炵懅閸樼數绱撻崒娆戝妽闁挎氨绱掑�???鍠氶悢鍡欐喐鎼粹埗鍝勵潨閳ь剚淇婇悽绋跨妞ゆ牭绲鹃弲婊堟⒑閸涘﹥澶勯柛�?�噹閳绘挾绱掑Ο鑲╃槇闂佽法鍣﹂敓锟?????閻庤娲栧ú銈夋偂閻斿吋鍊甸悷娆忓绾炬悂鏌涢弬鍧�?弰闁糕斁鍋撳銈嗗笒閸婂綊寮抽敓�?????濠电姷顣槐鏇㈠磻濡厧鍨濇繛鍡楁禋濞兼牜绱撴担鑲℃垶鍒婇幘顔界厽闁瑰浼濋鍕ㄦ灁閿燂�??閸曨兘鎷洪梺纭呭亹閸庢垿骞忛敓锟????闂佽法鍠嶇划娆撳箖瑜旈幃鈺呮嚒閵堝懐銈﹂梻濠庡亜濞诧妇绮欓幒�???鐤鹃柟闂寸劍閿燂�???? dcache 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮蹇涙偐缂佹ê娈ゅ銈嗗笒閸嬪棝宕�?ú顏呪拻濞达絽鎳欒ぐ鎺撴櫢闁跨噦锟?????濠碉紕鍋戦崐鎴﹀垂閻戞鈹嶆繛璇ф�??閿熻棄娲╅妵鎰板箳閹捐泛骞堥梻浣哥枃椤宕曢搹顐ゎ洸闁绘劦鍏涚换鍡涙煟閹板�?鎮嶉柟鍑ゆ嫹?闂佽法鍠撻弲顐﹀极椤旂晫�???闁告洦鍓﹂崑銊╂⒑閻愯棄鍔滈柡�?�偢�?�悂寮�?�?顒傛崲濠靛洨�???闁稿本绮岄敓�????闂備胶绮幐鍫曞磿閻㈢ǹ钃熼柨婵嗩槸閿燂拷??????????濠电姷鏁告慨鐑斤�??锟介鐐潟闁哄洢鍨圭壕濠氭煙鏉堝墽鐣辩痪鎯х秺閺岋拷?锟筋吋鎼达拷?锟界凹闂佸搫妫欑划宀勫煘閹达附鍋愰柛娆忣槸椤︹晠姊洪幖鐑囨嫹?閿熸枻锟???閿熸垝鍗冲璇测槈閵忊晜鏅濋梺鎸庣箓濡盯藝閵夆晜鈷戠紓浣股戠亸銊╂煕鐎ｎ偅宕屾慨濠勭帛閹峰懘宕ㄦ繝鍐ㄥ壍婵犵數鍋涢惇浼村垂閽樺鏆︾憸鐗堝笚閹偤鏌涜箛鎿冩Ц濞存粎鍋撻幈銊ヮ潨閸℃顫梺鎼烇�??锟藉ú锕傚箞閵婏妇�???闁告劏鏂傛禒銏狀渻閵堝啫鐏い銊ワ躬閺佹捇鏁撻敓�?????婵＄偑鍊栫敮鎺楀磹婵犳碍鍎楅柟鍓х帛閻撶喖鏌曡箛鏇炐ｉ柛鐔哄仱閺屾冻锟???閿熺瓔浜滈埀�???娼�?�濠氭晲婢跺﹥顥濋梺鍓茬厛閸犳宕愰鐐粹拺缂備焦蓱鐏忣厾绱掔紒妯哄闁糕晝鍋ら獮瀣晜閽樺姹楅梻浣藉亹閳峰牓宕滃☉銏╂晩濠电姴娲﹂埛鎴澝归崗鑲╂噮缂佸鍠栭湁婵犲﹤鍟伴崺锝忔�??閿熺瓔鍠栭�?�鐑藉极閹版澘閱囬柕蹇嬪灪濠㈡垿姊绘担鍛婃儓闁哥喓锟??瀹曟垿骞樼紒姗堟�??閿熶粙鐓崶銉ュ姢闁伙絿鏁婚弻鈥崇暆鐎ｎ偄锟???闂佽法鍠撻弲顐﹀汲閸℃稒鐓冪憸婊堝礈閻旈鏆�?ù鍏兼綑閿燂拷?????濠电姷鏁搁崑娑樜涘▎鎾冲瀭闁割偅娲栫粣妤呮煕閳╁啰鈯曢柣鎾寸懇閺岋綁骞嬮悘娲讳邯閹﹢鏁冮崒娑樹化闂佽婢樻晶搴ｅ鐠恒劎纾奸弶鍫涘妼濞搭喗銇勯�?锛勬噧闁宠閰ｉ獮鍡氼槼妞ゆ柨�?�板缁樻媴閸濄儲鐎┑鈽嗗亜鐎氭媽妫熷銈嗙墱閸庢垹绱為弽銊х瘈闂傚牊渚楅崕鎰版煛閸涱喚�???闁哄矉锟?????婵＄偑鍊戦崕鎻掔暆缁嬫娼栫紓浣股戞刊鎾煟閻旂厧浜伴柛銈咁儑缁辨挻鎷呯粵�?�闂佺ǹ锕ら�?�鐑藉箠閻愮儤鐒硷拷?锟姐儱妫�?▓鎰版⒑閸愬弶鎯堥悗姘煎墮閻剛绱撻崒姘炬嫹?閿熶粙宕愰悜鑺ワ�??锟介柨鏇氱缂嶆ê鈹戦悙鑼憼缂侇喖绉堕崚鎺戭吋婢跺á锕傛煕閺囥劌鐏犵紒鐘崇洴閺屽秵娼幏灞藉帯婵炲锟??缁犳牕顫忓ú顏呭仭闁哄�?�ч崐顖炴⒑閸涘﹥鈷愰柣鐔叉櫊閻涱喖螖閸涱參鍞堕梺鍝勬川閸嬫盯宕妸銉富闁靛牆妫欑亸鐢告煕閻樿櫕宕岋�??锟芥洏鍨介幐濠冨緞閸℃ɑ鏉告俊鐐�??锟介弻銊╋綖閺囩喓顩锋繝濠傜墛閻撴洟鎮楅敐搴′簼閻忓繑澹嗙槐鎺旂磼濡皷濮囬梺鐟板槻閹虫ê鐣烽敓锟???楠炴捇骞掑┑鍛；濠碉紕鍋戦崐鎰板疾閻樿缁╅弶鍫氭櫆�?�曞弶绻濋棃娑欏窛缂佲檧鍋撻梻浣呵归張顒傜矙閹存績鏋嶇憸蹇曟閹烘鍊锋い鎺嗗亾閿燂�??閸愵喗鐓曢悗锝庡亜婵淇婇崣澶婂妤犵偞顭囬埀顒佺⊕閿氭い搴㈡崌濮婅櫣鎷惔鈩冨劄鐟滅増甯掗惌妤呮煛閸ャ儱鐏柍閿嬪灴閺屾稖绠涢弴鐐蹭粯濡炪�?��?�╃划宥囨崲濞戞瑥绶為悗锝庡亞閿燂拷???濠碉紕鍋戦崐鏍暜婵犲嫭顐介柨鐔哄Т閻ゎ噣鐓崶銊р姇闁绘挻娲熼弻銊モ攽閸℃冻锟???閿熻姤绻涢崨顓犫枌闁瑰嚖�????闂佽法鍠曟慨銈吤洪敓�????瀹曞綊宕滄担鐟板簥濠电娀娼ч鍛存倷婵犲嫭鍠愰幖娣�?妽閸婂灚銇勯幒鎴濐仾闁抽攱鍨块弻锝夋偄閸涘﹦鍑￠梺鎶芥敱濮婅崵妲愰幒妤婃晪闁告侗鍘炬禒鎼佹�?�濞堝灝鏋熼柣鎿勭節閻涱噣寮介妸�???顎撻梺闈╁瘜閸樼厧顕ｉ幎鑺モ拻濞达綀娅ｇ敮娑欑箾閸欏澧碉拷?锟芥洩锟?????????
        .ren_o(backend_dcache_ren),
        .wstrb_o(backend_dcache_wen),
        .writen_o(backend_dcache_writen),
        .llw_to_dcache(llw_to_dcache),
        .scw_to_dcache(scw_to_dcache),

        .virtual_addr_o(backend_dcache_addr),
        .wdata_o(backend_dcache_write_data),

        .is_exception_execute1(is_exception_execute1),
        .rdata_i(dcache_rdata),
        .rdata_valid_i(dcache_backend_rdata_valid),
        .sc_cancel_to_backend(sc_cancel_to_backend),
        .uncache_i(uncache_out),
        .dcache_pause_i(~dcache_ready),
        .dcache_is_exception_i(dcache_is_exception),
        .dcache_exception_cause_i(dcache_exception_cause),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸パ勶拷?锟介悗骞垮劚閹峰宕ワ拷?锟筋喗鐓曢柍鈺佸暞锟??鍫㈢磼閻樺啿鍝烘慨濠冩そ瀹曘劍绻濋崟�???娅戞俊鐐拷?锟斤�??锟藉矂宕归柆宥呯疄闁靛ǹ鍎洪崥瀣煕閿燂拷?閺呮粓顢欓弮鍫熲拺缂備焦锚婵牊绻涢崗鑲╂噧闂囧鏌ㄩ悤鍌涘�???濠电偛鐗嗛悘婵嗏枍閿燂拷?閺屾盯骞樼捄鐑樼亪濡ょ姷鍋涢崯顐�?煝鎼淬劌绠奸柛鎰ㄦ櫆濞呭矂姊婚敓�????閳ь剛鍋涢懟顖涙櫠椤栫偞鐓曢柟鐑樺�?闊剚顨ラ悙鑼фい銏＄懇瀹曟粏顧傜紒杈ㄥ▕濮婄粯鎷呴崨闈涚秺瀵敻顢楅崟�???浠悷婊勬煥閻ｅ嘲鈹戦崱鈺佹倯闂佹悶鍎弲婵嬫晬濠婂牊鐓熼幖鎼灣缁夌敻鏌涳�??锟筋亜顏柟顔筋焽閳ь剚绋掕彠濞存粍绮撻弻鏇＄�?閵壯咃紵婵犫拃鍜佹殰闁瑰嚖锟???闂佽法鍠曟慨銈吤哄Ο鍏兼殰闁跨喓濮寸粻鏍ㄧ箾閸℃ɑ灏伴柛銈嗗灦閵囧嫰骞掗幋顖氬濡ょ姷鍋戦崹钘夘潖婵犳艾纾兼繛鍡樺姉閵堟澘顪冮妶搴�?�簻妞わ富鍨堕弫鎾绘晸閿燂拷????婵＄偑鍊戦崹鐑樼┍濞诧拷?锟藉洩銇愰幒鎾跺幍濡炪�?�姊归崕铏闁�?秵鐓欐い鏃囧吹閻瑱�????閿熻姤娲忛崝宥囨崲濠靛�?嬫い鎰╁灮椤�?垿姊婚崒姘炬�??閿熶粙鎳楅崜浣稿灊妞ゆ牗鍑瑰鏍棯椤撶偞鍣峰ù婊冪秺閺屾盯骞囬妸锔界彇濡炪�?�鏅炵亸娆戞閹烘梹宕夐柣鎴灻弸鐘测攽椤旂》宸ユい顓炲槻閻ｇ兘骞掗幋顓熷兊濡炪倖鍨煎Λ鍕妤ｅ啯鐓欓梻鍌氼嚟椤︼妇鐥幆褏绉洪柡锟??鍠栧浼欐嫹?閿熻棄澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鎴﹀箰閹惰棄钃熼柨娑樺濞岊亪鏌涢幘妞诲亾婵℃彃鐗撳鐚存嫹?閿熺晫濯鎰版煕閵娿儳浠㈤柣锝囧厴瀹曪繝鎮欏鍡樷拹缂佺粯绻冮幏鍛存惞閻у摜闂梻鍌氾拷?锟介崐宄懊归崶顒夋晪鐟滄繈骞忛敓�?????闂佽法鍠曡闁哄懏鐩敐鐐测攽鐎ｏ拷?锟解晠鏌ㄩ弮鍥撻柣婵嗗槻閳规垶骞婇柛濠冩礋楠炲﹥鎯旈姀鈺傛暞闂傚�?�鍊风粈�???骞夐垾瓒佹椽鏁冮崒姘拷?锟介梻渚囧墮缁夋挳鎮块悙顒傜瘈濠电姴鍊绘晶娑㈡煕鐎ｅ墎绉�?柡灞剧洴婵＄兘顢欓懡銈囨晨闂備焦鐪归崝宀勫箹椤愶附绠掗梻浣虹帛鏋繛鍛礈娴滄悂鏁傞懞銉ュ伎婵犵數濮撮幊蹇涱敂閻樼粯鐓欏�?�閳诲牓鏌熷畷鍥р枅妞ゃ垺顨婂畷鎺�?Χ閸涱喗姣嗗┑鐘殿暜缁辨洟宕戦幋锟??纾归柡宥庡幖閸ㄥ倿鏌ｉ姀鈩冪秳闁搞儺鍓﹂弫宥夋煟閹存繃宸濈紒瀣箻濡懘顢曢�?鈥愁槱闂佺懓鍢查鍛弲濡炪倕绻愮粔鐢稿疾濠婂牊鈷戦柛娑橈攻婢跺嫬霉濠婂懎浠遍柟顔界懄缁绘繈宕堕妸銏″濠电偠鎻徊浠嬪箟閿熺姴鐤柣鎰嚟缁犻箖鎮归崶鍥ф噽閺嗐倝鎮楃憴鍕闁搞劌鐏濋悾鐑藉Ω閳哄﹥鏅ｅ┑鐐村灦閻熝勭閺嶃劋绻嗛柣鎰典簻閳ь剚鐗犻獮鎰板醇閺囩偛鐎┑鐐叉▕娴滄粓鎮￠弴銏＄厵閻庣數枪鍟哥紒鐐礃濡嫰�?�?梺鎸庣箓濞诧箓顢旈悢鍑ゆ�??閿熻棄顫濋鐘缂備胶绮惄顖氱暦婵傚憡鍋勯柛鎾冲级椤ュ牓姊绘担鍛婃儓閻炴凹鍋婂畷婵嬪箣濠垫劕娈ㄩ梺鍦檸閸犳牗鍎梻�???娼ч悧鍡椕洪妸銉㈡灃闁秆勵殕閳锋帒霉閿濆妫戝☉鎾瑰皺缁辨帡骞撻幒鎾充淮闂佽法鍣﹂敓锟??????闂佽法鍣﹂敓�?????????婵＄偑鍊栧Λ浣肝涢崟顒傤洸闁荤喖鍋婂�?�濠氭煏閸繃顥滃┑顕嗙畵閺佹捇鏁撻敓锟?????婵犵數濮伴崹濂革綖婢跺⊕娲偄婵傚缍庡┑鐐叉▕娴滄粎绮绘导鏉戠閺夊牆澧介幃濂告煟閿濆懐浠涘ǎ鍥э躬婵″爼宕堕‖顔哄灲閺岀喓鎷犺绾捐法绱掗纰卞剰妞ゆ挸鍚嬪鍕舵嫹?閿燂�??锟藉煐閿燂拷??闂佽法鍠嶇划娆撳蓟閿濆顫呴柕蹇婂墲濮ｅ嫰姊洪幐搴ｂ姇缂侇喗鎸搁～蹇涙惞閸︻厾锟????闂佽姘﹂～澶娒哄⿰鍫濇瀬濠电姵鑹剧粻鏍煙椤栵絿浜规繛宸憾閺佸�?�鏌涘☉鍗炵仩妤犵儑�??????闂備緤锟???閿熻棄鑻晶鎾煥閻曞�?�锟???婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓熷濠氼敍閻愬鍙嗛梺鍝勬川閸庢垿骞忛敓�?????闂佽法鍠撻弲顐ゅ垝婵犳凹鏁嶉柣鎰嚟閸欏棝鏌ㄩ悤鍌涘�??????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犲灚鍔栧瓭闂備緤�????閿熻棄鑻晶鍓х磼閻樿櫕灏柣锝囧厴�?�曞ジ寮撮妸锔芥珜闂備緤�????閿熻棄鑻晶鎵磼椤旂⒈鐓奸柟顔规櫇缁辨帒螣閻撳骸绠為梻鍌欑窔閳ь剚绋戝畵鍡樼箾娴ｅ啿娲ら崙鐘绘煟閺傚灝鎮戦柣鎾跺枛閺�?喖骞戦幇顓狅�??锟介梺鍝勵儐閻╊垶寮婚敐澶婄闁告劑鍔嬮崰濠囨�?�鐟欏嫭�?夐柛鈺傜墵钘濋柣�???鐗婇崕鐔兼煃閽樺顥滄繛鍫濄偢濮婂宕掑顑藉亾妞嬪孩顐介柨鐔哄Т閻骞栧ǎ锟??濡奸柛銊ワ拷?锟介弻娑㈩敃閿濆棛顦ラ梺钘夊暟閸犳牠寮诲澶娢ㄩ柕澹秶�?婇梻浣告惈濡螞濠靛绠栨俊銈呮噺閺呮煡骞栫划鍏夊亾閹颁焦楠勯梻鍌欐缁鳖喚绮婚幋锔藉亱闁规崘顕х粻鏍ㄤ繆閵堝懎鏆為柛鐘叉閺屾盯寮撮妸銉ヮ潾闂佹寧绋掗敃銏�?潖濞差亜宸濆┑鐘插暊閹峰綊姊洪幖鐐插婵炲皷鍓濇穱濠忔嫹?閿熻姤蓱婵绱掗娑欑闁诲骸顭峰娲捶椤撶偘澹曞┑鐐插悑閻熲晠骞嗛崒鐐茬妞ゆ帒鍊婚惁鍫ユ⒑闂堟盯鐛滅紒鎻掑⒔濞戠敻鎮欓璺ㄧ畾濡炪�?�鍔х紞鍡椻枔閺囩姷纾奸柛灞炬皑鏍￠梺闈涚墳缂嶄礁鐣烽敓锟???閸╋繝宕�?妸銉ь吋闂傚�?�鍊峰ù鍥綖婢舵劦鏁婇柡宥庡幖缁愭鏌�?�搴�?�伎闁瑰嚖锟???闂佽法鍠曟慨銈囩紦娴犲宸濆┑鐘插楠炴姊绘担绛嬫綈闁稿孩濞婇、姘额敇閻忕粯妞介獮�???顢欓悾灞藉箥婵＄偑鍊栧褰掑几婵犳碍�???闁秆勵殕閻撴瑦銇勯弮鍌涙珪闁瑰啿瀚伴弻銊モ槈濞嗗繐顫岄梺瀹狀潐閸ㄥ灝鐣烽崡鐑嗘建闁糕剝顨嗛弳銏＄�?閻㈤潧啸闁轰礁鎲￠幈銊╂偨閸撳弶鏅╅梺鍝勭▉閸樿偐绮ｅΔ鍛厸鐎广儱楠搁獮鏍棯閹呯Ш闁哄本绋栭ˇ铏亜閵娿儲鍤囬柟閿嬪灴閹垽宕楅懖鈺佸箺闂備礁鎼崯顐﹀磹閻㈢ǹ绠柨鐔哄У閻撴稑霉閿濆浜ら棅顒夊墴閺岋拷?锟界暆鐎ｎ剙鍩屽銈庡亝缁诲牓銆佸Δ鍛＜婵炴垶鐟ラ弸娑㈡⒒娴ｇ瓔鍤欓悗娑掓櫊閺佹捇鏁撻敓�????????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏缂佸鍨剁粋鎺撶附閸涘ň鎷虹紓鍌欑劍閿氶柣蹇氶哺娣囧﹪顢曢姀�???�???缂備緡鍠栭�?�鐑界嵁鎼淬劍鍤嶉柕澹啫绠ラ梻浣筋嚙鐎涒晝绮欓幒鏇熸噷闂備焦濞婇弨閬嶅礉閺嶎厼桅闁告洦鍨奸弫鍐煏韫囧﹥鍤曢柕蹇嬶�??锟介悡鍐偡濞嗗繐顏╅柣蹇撶摠閵囧嫰�???閿涘嫭鍣紓渚囧枤椤ｎ噣骞忛敓锟????闂佽法鍠撻悺鏃堝磻閸℃稑姹查柕澶涘閿燂�??缂佸墽澧楄摫妞ゎ偄锕弻娑虫�??閿熺瓔浜濋崳褰掓懚閻愮儤鐓曢柟浼存涧閺嬫盯鏌★拷?锟解晝绐旈柡�???鍠栧畷婊嗩槾閻㈩垱鐩弻锟犲川椤�?枻锟???閿熶粙鏌＄仦璇插闁诡喓鍊濆畷鎺戔槈濮楀棔锟???8濠电姷鏁告慨鐑藉极閸涘﹥鍙忛柣鎴ｆ閺嬩線鏌涘☉姗堟敾闁告瑥绻橀弻锝夊箣閿濆棭妫勯梺鍝勵儎缁舵岸寮诲☉妯锋婵鐗婇弫楣冩⒑閸涘﹦鎳冪紒缁橈�?��?�鏁愭径濠勵吅闂佹寧绻傚Λ顓炍涢崟顖涒拺闁告繂瀚烽崕搴ｇ磼閼搁潧鍝猴拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝棎浜滄い鎾跺Т閸樿揪�????閿熺瓔鍠栭�?�鐑藉极閹版澘宸濋柛灞剧矊閺嬪酣鏌嶇拠鏌ュ弰妤犵偛妫滈ˇ铏亜閺傚灝顏紒杈ㄦ崌�?�曟帒鈻庨幒鎴濆腐濠电姵顔栭崰妤呭箰閹惰棄绠栨俊顖欒濞尖晠鎮规潪鎵Э闁挎洖鍊归悡鏇㈡煛閸ャ儱濡奸柡瀣舵�???闂傚倸鍊风粈浣革耿闁�?秴纾婚柟鎹愵嚙缁犳岸鎮橀悙璺衡枏婵炴垯鍨洪崐鐑芥煟閵忋垺鏆╅柨娑欑箖缁绘稒娼忛崜褎鍋ч梺鍝勬媼閸嬪﹤鐣锋總鍓叉晜闁割偆鍠撻崢杈ㄧ節閻㈤潧孝闁哥喐澹嗙划濠氭倻閸ャ劌�????闂佽法鍠撻悺鏃堝窗閺嶎叏�????閿熶粙鎮滈挊澶嬶�??锟介梺褰掑亰閸樿偐娆㈤悙鐑橈�??锟介柨婵嗛�?�娴滄繈鏌ｅ┑鍥р枙婵﹦绮幏鍛村川婵犲倹娈樺┑鐐存尰绾板秹銆冩繝鍌滄殾鐟滅増甯楅幆鐐淬亜閹扳晛鐒洪柛銈冿拷?锟藉娲箹閻愭彃濮堕梺鍛婃尰锟??鎼佸春濞戙垹绠ｉ柣鎰暩椤旀洟姊洪悡搴涘仮妞ゃ�?�鍊垮畷闈涒枎閹板灚顔旈梺缁樺姈閹苯鈻撳⿰鍫熺厸閿燂拷?閳ь剟宕伴弽顓犲祦闁哄秲鍔嶆刊鎾煣韫囨凹娼愭慨锝呮处娣囧﹪濡堕崶顬儵鏌涳拷?锟筋偆娲撮挊婵嬫煟閵忕姵鎲革�??锟芥挷绶氶弻鈥愁吋閸愩劌顬夋繝娈垮灡閹告娊寮婚敐澶嬪亜缁炬媽椴稿▓銉х磽閸屾艾鏆炴繛鑼�?枎椤繒绱掑Ο璇诧�??锟界紓浣割儐椤戞瑥螞�???鍕拺缂佸顑欓崕蹇涙煙閾忣偄濮嶆鐐村灴閿燂拷?闁靛牆鎳愰ˇ鏉款渻閵堝棛澧紒瀣灦缁傛帡顢橀�?�???鎷洪梻鍌氱墛閸楁洟宕奸妷銉ф煣濠电姴锕ら悧鍡涙偂閺囥垺鐓欓弶鍫ョ畺濡绢噣鏌ｉ幘瀛樼缂佺粯绻堝Λ鍐ㄢ槈濞嗘ɑ顥ｆ俊鐐�??锟界换鎴�?箰閹惰棄钃熸繛鎴炵懄閸庣喖鏌嶉埡浣告殲鐎规洖纾槐鎾存媴娴犲鎽甸柣銏╁灲缁绘繈鐛繝鍌�?牚闁割偆鍣ュΛ鍐ㄢ攽閻愭潙鐏﹂拑閬嶆煙閾忣偆鎳囬柡�?嬬稻閹棃锟??閳轰焦娅涢梻浣告憸婵敻鎮ч悩璇茬伋闁挎洖鍊归崐濠氭煢濡警妲洪柣锝嗘そ濮婃椽妫冨☉姘辩杽闂佺ǹ锕ラ悧鐘茬暦閹达箑纾奸柣鎰皺椤�?劙鏌℃径濠勫濠�?呮櫕缁棃鎮介崨濠勫幈闂佺粯鍔樼亸娆戠矓閻戞ɑ鍙忓┑鐘插鐢稓绱掑Δ鍐ㄦ灈闁糕斁鍋撳銈嗗笒鐎氼剟鎮為崹顐犱簻闁瑰搫绉烽崗�?勬煃閽樺妾ч柟鍑ゆ嫹?闂佽法鍠曟慨銈夊箰缁嬭娑樷枎閹寸偛搴婂┑鐐村灦閻燂附鍒婇幘顔界厱闁归偊鍘肩徊濠氭煛閸℃韬柡�?嬬磿閳ь剨缍嗛崑鍛村煕閹扮増鐓忛柛銉戝喚浼冨Δ鐘靛仦椤洭骞戦崟顒佸闁绘鐗忓鏍⒒閸屾瑦绁伴柕鍡忓亾闂佺ǹ顑嗛幐鎼佹箒闂佺粯锚濡﹪宕曢幇鐗堢厽闁规儳鍟块弳锝夋煛锟??瀣暠閾伙絽銆掑鐓庣仭閺佸牊淇婇悙顏庢�??閿熶粙宕曢懠�???鍨濋敓锟???閸曨剛鐣冲┑鐘垫暩婵挳鏁冮妶鍥ｅ亾濮樼厧鏋ょ紒顔碱煼閹瑩鎮滃Ο鐓庡箰闂佽绻掗崑鐘活敋瑜庨幈銊╁磼閿旇棄锟???闂佽法鍠撻悺鏃堝窗閿燂拷?椤洤鈻庨幒鏂捐埅闂佽法鍣﹂敓锟????????缂傚倷娴囨ご鎼佹偡閳哄懎钃熼柨婵嗘閸庣喖鏌曡箛濠冩珔闁哄懘浜跺娲传閵夈儛锝夋煥閻曞倹锟??????闂佽娴烽幊鎿勬�??閿熸垝鍗冲畷鎴炵�?閸パ冩優闂佸搫娲㈤崹娲偂濞嗘垹纾藉ù锝夋涧閻忊晠鏌★�??锟筋偆鈯曢柕鍥у椤㈡洟锟??閳ヨ櫕鐣婚梻浣告惈閻寰婇崐鐔轰航婵犵數鍋涘Λ娆撳磿閸愭祴鏋�?い鎾卞灪閳锋垿寮堕悙闈涱暭缂佷胶澧楅妵鍕敃閵忊晜楔闂佺懓绠嶉崹褰掑煘閹寸姭鍋撻敐搴′簻濞寸姵妞藉濠氬磼濮樺崬�???缂備礁顑呴悧鎾愁嚕閹间礁宸濇い鎾寸⊕閿燂�??闂備胶绮崝鏍ь熆濡棿鐒婇柛鎰靛枟閻撴洟鐓崶銊︾鐎涙繄绱撻崒姘毙㈤柨鏇橈�??锟介幃楣冩�?�閽樺顔婇梺鐟扮枃閸╂牜鏁�?垾宕囨殾婵°�?�鎳忛崵鍐煃閸濆嫸�????閿熶粙宕归柆宥嗏拻濞达絿鐡旈崵鍐煕閻樻剚娈滈柟顔惧厴閸╋繝宕ㄩ鐘垫毇婵犵數濮撮敃銈夊触閿燂拷?閹垽宕楅懖鈺佸汲闂佽鍑界紞鍡樼閼搁潧顕遍柡宥庡幗閳锋帡鏌涚仦鍓ф噭缂佷焦澹嗛�?顒冾潐濞叉牠鎮樺璺虹疄闁靛ň鏅涢崹鍌涖亜閹扳晪锟???閿熻棄煤閸涘﹦绠鹃悗鐢登瑰瓭濡炪倖鍨甸幊鎰垝閸喎绶為柟閭�?幖閳ь剙鐖奸弻锝夊箛椤斿墽顦伴梺鍦劋椤ㄥ懘宕欓悩纰樺亾楠炲灝鍔氭い锔垮嵆閹�??锟解枎閹惧鍘靛┑鐐茬墕閻忔繈寮稿☉娆嶄簻闁挎繂鎳岄崑銏ゆ煛�???瀣М妤犵偞顭囬埀顒勬涧閹诧繝宕虫导�?�樷拺闁告繂瀚﹢浼存煟閳哄﹤鐏﹂柣娑卞枤閳ь剨缍嗘禍鏍几鎼淬劎鍙撻柛銉戝秴浼愭繛�?�樼矒缁犳牠寮婚垾鎰佸悑閹艰揪锟???閿熺晫鐖遍梻浣呵归鍡涘箰閹间緤缍栨繝闈涱儐閿燂�??????
        .flush_o(flush_o),
        .pause_o(pause_o),

        .icacop_en(icacop_en),
        .dcacop_en(dcacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),
        
        //debug
        .debug_wb_valid1(debug_wb_valid1),
        .debug_wb_valid2(debug_wb_valid2),
        .debug_pc1(debug_pc1),
        .debug_pc2(debug_pc2),
        .debug_inst1(debug_inst1),
        .debug_inst2(debug_inst2),
        .debug_reg_addr1(debug_reg_addr1),
        .debug_reg_addr2(debug_reg_addr2),
        .debug_wdata1(debug_wdata1),
        .debug_wdata2(debug_wdata2),
        .debug_wb_we1(debug_wb_we1),
        .debug_wb_we2(debug_wb_we2) 


        // difftest
        `ifdef DIFF
        ,

        .diff0              (diff0              ),
        .diff1              (diff1              ),
        .stable_counter     (cnt                ),

        .regs_diff          (regs_diff_out      ),

        .csr_crmd_diff      (csr_crmd_diff_0    ),
        .csr_prmd_diff      (csr_prmd_diff_0    ),
        .csr_ectl_diff      (csr_ectl_diff_0    ),
        .csr_estat_diff     (csr_estat_diff_0   ),
        .csr_era_diff       (csr_era_diff_0     ),
        .csr_badv_diff      (csr_badv_diff_0    ),
        .csr_eentry_diff    (csr_eentry_diff_0  ),
        .csr_tlbidx_diff    (csr_tlbidx_diff_0  ),
        .csr_tlbehi_diff    (csr_tlbehi_diff_0  ),
        .csr_tlbelo0_diff   (csr_tlbelo0_diff_0 ),
        .csr_tlbelo1_diff   (csr_tlbelo1_diff_0 ),
        .csr_asid_diff      (csr_asid_diff_0    ),
        .csr_save0_diff     (csr_save0_diff_0   ),
        .csr_save1_diff     (csr_save1_diff_0   ),
        .csr_save2_diff     (csr_save2_diff_0   ),
        .csr_save3_diff     (csr_save3_diff_0   ),
        .csr_tid_diff       (csr_tid_diff_0     ),
        .csr_tcfg_diff      (csr_tcfg_diff_0    ),
        .csr_tval_diff      (csr_tval_diff_0    ),
        .csr_ticlr_diff     (csr_ticlr_diff_0   ),
        .csr_llbctl_diff    (csr_llbctl_diff_0  ),
        .csr_tlbrentry_diff (csr_tlbrentry_diff_0),
        .csr_dmw0_diff      (csr_dmw0_diff_0    ),
        .csr_dmw1_diff      (csr_dmw1_diff_0    ),
        .csr_pgdl_diff      (csr_pgdl_diff_0    ),
        .csr_pgdh_diff      (csr_pgdh_diff_0    )
        `endif      
    );

    wire icache_ren_received;
    wire dcache_ren_received;
    wire icache_flush_flag_valid;

    wire iuncache_rvalid;
    wire [63:0] iuncache_rdata;
    wire iuncache_ren;
    wire [31:0] iuncache_raddr;

    wire [31:0] inst_paddr;
    wire iuncache_en;

    wire inst_addr_trans_en;
    icache u_icache
    (
        .clk(aclk),
        .rst(rst),   
        .flush(flush_o[1]),       
    // Interface to CPU
        .inst_rreq(inst_rreq),  
        .not_same_page(not_same_page),
        .iuncache_en(iuncache_en),
        .inst_addr1(inst_addr1),   
        .inst_addr2(inst_addr2),  
        .paddr(inst_paddr),
        .if_pred_addr1(if_pred_addr1),
        .if_pred_addr2(if_pred_addr2),
        .BPU_pred_taken(BPU_pred_taken),

        .icacop_en(icacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),

        .pi_is_exception(pi_is_exception),
        .pi_exception_cause(pi_exception_cause),
        .inst_addr_trans_en(inst_addr_trans_en),
        .inst_tlb_found(inst_tlb_found),
        .inst_tlb_v(inst_tlb_v),
        .inst_tlb_plv(inst_tlb_plv),
        .csr_plv(csr_plv), 

        .pred_addr1(pred_addr1_for_buffer),
        .pred_addr2(pred_addr2_for_buffer),
        .pred_taken(pred_taken_for_buffer),
        .inst_valid1(icache_inst_valid1),  
        .inst_valid2(icache_inst_valid2),   
        .inst_out1(icache_inst1),       
        .inst_out2(icache_inst2),
        .valid_out(icache_valid_out),
        .pc1(icache_pc1),
        .pc2(icache_pc2),
        .pc_is_exception_out1(pi_icache_is_exception1),
        .pc_is_exception_out2(pi_icache_is_exception2), 
        .pc_exception_cause_out1(pi_icache_exception_cause1),
        .pc_exception_cause_out2(pi_icache_exception_cause2),
        .pc_suspend(pc_suspend), 
    // Interface to Read Bus
        .dev_rrdy(dev_rrdy_to_cache),       
        .cpu_ren(icache_ren),       
        .cpu_raddr(icache_araddr),      
        .dev_rvalid(icache_rvalid),     
        .dev_rdata(icache_rdata),
        .ren_received(icache_ren_received),
        .flush_flag_valid(icache_flush_flag_valid),

        .uncache_rvalid(iuncache_rvalid),
        .uncache_rdata(iuncache_rdata),
        .uncache_ren(iuncache_ren),
        .uncache_raddr(iuncache_raddr)   
    );

    wire debug_wb_valid1;
    wire debug_wb_valid2;
    wire [31:0] debug_pc1;
    wire [31:0] debug_pc2;
    wire [31:0] debug_inst1;
    wire [31:0] debug_inst2;
    wire [4:0] debug_reg_addr1;
    wire [4:0] debug_reg_addr2;
    wire [31:0] debug_wdata1;
    wire [31:0] debug_wdata2;
    wire debug_wb_we1;
    wire debug_wb_we2;

    wire [3:0] duncache_wstrb;

    wire cache_axi_write_pre_ready;
    wire duncache_en;
    wire data_fetch;

    wire data_addr_trans_en;
    dcache u_dcache(
        .clk(aclk),
        .rst(rst),
        .bvalid(bvalid),
        
        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓顕崑娑⑺夊鑸电厱婵炲棗绻戦幆鍫ユ煃鐟欏嫬鐏撮柟顔规櫊瀹曞綊顢曢敐鍡欐婵犵數濮甸鏍窗濮樿泛绀傛慨妞诲亾濠碘剝鎸冲畷鎺戔槈濮樺吋绁梺璇插嚱缂嶅棙绂嶉悙鏍稿洭顢橀悙鈺傛杸闂佺粯顭囩划顖氣槈瑜庨妵鍕箣濠靛洤娅х紓渚囧枛椤嘲顕ｆ禒�?�垫晣闁绘柨鎼獮鍫ユ⒑鐠囪尙绠抽柛瀣⊕閺呰埖绂掞�??锟筋亞鍘介梺闈涳紡閸涱垽绱查梺鑽ゅТ濞层�?�顕ｉ崼�???澶愬閵堝棛鍘搁悗鍏夊亾閻庯綆鍓涜ⅵ婵°�?�濮烽崑娑㈩敄婢舵劕鏋侀柟鐗堟緲瀹告繈鏌涘☉鍗炴灍鐎规洖鐭傞弻鈥崇暆鐎ｎ剛鐦堥悗瑙勬磸閸�?垿銆佸▎鎾崇鐟滃繘宕㈤幒鏃傜＝闁稿本鐟︾粊鏉款渻鐎涙ɑ鍊愭鐐村姈缁绘繂顫濋鍌ゅ數闂備礁鎲＄粙鎴︽偤閵娾晛纾块敓锟???閳ь剛妲愰幒鏂哄亾閿濆簼绨藉ù鐘灮閹叉悂寮堕幐搴闂佸疇顫夐崹鍫曠嵁婵犲洦鐓曞┑鐘插枤濞堟洟鏌熸鏍帨闁瑰嚖锟???闂佽法鍠曞Λ鍕箟閳ュ磭鏆﹂柛娆忣槷缁诲棙銇勯弽銊ф噯妞ゆ帞鍠愮换娑㈠礂閼测晛鈷堢紓浣介哺閹稿骞忛崨�?�樺殐闁斥晛鍟悘锕傛煕閹烘垟搴烽柟鍑ゆ�??闂佽法鍠曞Λ鍕箺濠婂懎顥氶柛蹇氬亹缁犻箖鏌燂�??锟界ǹ鍓冲〒姘洴閺屾稒鎯旈敍鍕唹缂備胶绮惄顖氱暦婵傚壊鏁冮柕蹇曞Х椤旀帞绱撻崒娆愮グ濡炲瓨鎮傞獮鎰節濮橆剛顔嗛梺鍛婄☉閻°劑骞嗛悙鐑樼厽闁绘梻枪椤ュ銇勯幇顑惧仮婵﹦绮幏鍛村川婵犲�?�娈樻繝娈垮枛閿曘�?�绱炴繝鍥ラ柛鎰ㄦ櫇閿燂拷?闂佹悶鍎�?弲娑氱矈閿曞倹鈷戠痪顓炴噺瑜把呯磼閻樺啿鐏撮柨婵堝仱瀹曨煉锟???閿熻姤顭囬崢顏堟⒑閸撴彃浜濈紒璇插暣瀹曠敻宕堕浣哄幈闂佺粯鍔樼亸娆撳春閿濆棙鍙忓┑鐘插暞閵囨繃淇婇銏犳殭闁宠棄顦板蹇涘Ω閹扳晪锟???閿熻棄顫忛搹鍦煓闁割煈鍣崝澶嬬節閻㈤潧浠滈柨鏇樺妼铻為柣鏂款殠濞撳鏌曢崼婵囶棡缁惧墽鏁婚弻娑虫�??閿熺瓔鍋呯亸浼存煙娓氬灝濡界紒缁樼箞瀹曘劑顢氶崨�???鎽嬪┑鐘垫暩閸嬬偤宕硅ぐ鎺戞瀬閻犲洩灏欓弳锕傛煏婵炵偓娅撻柡浣革躬閺屾稖绠涢幘鍗炰划闂佽桨绶℃禍婵堟崲濠靛鍋ㄩ梻鍫熷垁閵夛负浜滈柨婵嗗閻瑩鏌ㄩ悤鍌涘?婵＄偑鍊栫敮鎺楀疮椤栫偞鍋熸い蹇撶墛閻撴瑩鏌涜箛鏇炲付濠殿喖绉归弻鈥崇暆鐎ｎ剛袦闂佽桨鐒﹂崝娆忕暦閸洖惟闁挎梻鏅Σ妤呮⒒閸屾瑦绁版俊妞煎姂閹偤鏁冮崒姘鳖唹闂佹悶鍎洪崜娆撳几閿燂�??閺岀喖宕滆鐢盯鏌￠崨顔斤�??锟介柡宀嬫嫹???闂傚倸鍊搁崐鎼佸磹閻戣姤鍤勯柛鎾茬閸ㄦ繃銇勯弽顐粶缂佺姴缍婇弻宥夊传閸曨剙娅ｇ紒鐐礃椤曆囧煘閹达附鍋愰悹鍥囧嫬�????闂佽法鍠嶇划娆忣嚕閹惰姤鏅濋柛灞剧�?�閸樺崬顪冮妶鍡�?Ё缂佹煡绠栭弫鎾绘晸閿燂拷??闂備浇顕栭崹鎶藉窗閺嶎厼绠栵�??锟藉嫭澹嬮崼顏堟煕閹邦喖浜鹃弫鍫ユ⒒閿燂�??閳ь剚绋撻埞鎺楁煕閿燂�??閸ㄧ敻鎮鹃悜钘夐唶闁哄洢鍔嶉弲銏＄箾鏉堝墽鍒帮拷?锟筋喖澧庨埀顒佷亢閸嬫劗妲愰幘璇茬＜婵炲棙鍩堝Σ顔碱渻閵堝棗鐏ユ俊顐ｇ箞閵嗕線寮�?�閺嬪酣鏌熼幆褏锛嶉柨娑氬枎閳规垿鎮欓弶鎴犱桓闂佸磭顑曢崐婵嬪箖閿燂拷???闂傚倷绀�?幉鈥趁洪敃鍌氬偍濡わ絽鍟崑顏堟煕閺囥劌澧扮紒锟??鍋撶紓浣哄亾濠㈡﹢藝鏉堚晛顥氶柛褎顨嗛悡娑樏归敐鍥╂憘闁搞�?�鐟╅弻锝夋晲閸パ冨箣闂佽鍠撻崹濠氬窗婵犲啯缍囬柕濠忛檮閻濐偄鈹戦悩鎰佸晱闁哥姵顨婇弫鍐煛閸涱厾顦┑鐐叉閹告悂寮搁敓�????閺屾洟宕煎┑鎰ч梺鎶芥敱鐢帡婀�?梺鎸庣箓閹冲繒鎷归敓鐘虫櫢闁跨噦�????婵炲濮撮鍡涙偂閺囥垺鐓忓┑鐐茬仢婵¤姤銇勯妷銉Ч闁靛洤瀚伴、锟??鎮欙�??锟界硶鏁嶉梺璺ㄥ櫐閿燂拷??????闂備礁鎼ú鐘诲礈濠靛鏁傞柣妯款梿瑜版帗鍋戦柛娑卞弾濞差參姊洪悷鏉跨骇闁瑰憡濞婂顐�?箛閺夊灝鑰垮┑鈽嗗灣缁垳娆㈤锔解拻闁稿本鑹鹃�?顒傚厴閹虫宕滄担绋跨亰濡炪倖鐗滈崑娑氱矆婢跺绻嗘い鏍仦閿涚喖鏌ｉ幒鎴敾缂佺粯鐩畷鍗炍熼崫鍕垫綌婵犵數鍋涢幊鎰箾閳ь剚鎱ㄦ繝鍐┿仢妞ゎ澁�????缂傚倷绀�?ˇ閬嶅极婵犳艾绠栭柨鐔哄Т閸楁娊鏌曡箛銉х？闁告﹩浜濈换婵嬫偨闂堟稐绮堕梺璇茬箲缁诲啯绌辨繝鍥ㄥ仼閿燂�??閳ь剙螞椤栨稏浜滈柟鎹愭硾瀛濇繛�?�樼矒缁犳牠寮婚弴銏犵�?�鐟滃秹顢旈鐔翠簻闁靛繆鍓濈粈瀣煥閻曞�?�锟???闂備線娼х换鍫ュ春閸曨垰鑸归柧蹇撴贡绾句粙鏌涚仦鍓ф噭缂佷焦婢橀—鍐级閹寸偞鍠愰梺杞扮贰閸ｏ綁鐛幒锟??鍗抽柣妯跨簿閸╁懘姊婚崒娆愮グ鐎规洖鐏氶幈銊╁级閹炽劍妞芥俊鍫曞川閸屾粌鏋戠紒缁樼箞瀹曟儼顦撮柛鏃撶畱椤啴濡堕崱妤冪憪闂佺粯甯粻鎴︽偩妞嬪簼娌柣鎰靛墮瀵寧绻濋悽闈浶㈤柛鐕佸灦婵￠潧鈹戦幘鏉戭伓?闂佽法鍠曟慨銈吤洪敓�????閵嗗啯绻濋崒銈嗙稁闂佺厧顫曢崐鏇⑺夊鑸碉拷?锟介柨婵嗙凹缁ㄤ粙鏌涢弮鍌涙毈婵﹤顭峰畷鎺戔枎閹烘垵锟???闂備浇顕э�??锟解晝绮欓崼銉ョ柧婵犲﹤鎳忓畷鍙夌箾閹寸偟鎳呯紒�???鍋撻梻浣告啞閸擃剟宕ㄩ婊勬瘞闂傚�?�娴囬褝锟???閿熻В鏅濈划娆撳箳濡炵儵鍋撻敃鍌氱倞闁宠桨�?佽ⅲ闂備緤锟???閿熻棄鑻晶瀛樻叏婵犲啯銇濇鐐寸墵閹瑩骞撻幒鎴綑闂傚�?�绀�?幉锟犲蓟閵娾敡鍥偨閸濄儱绁﹂棅顐㈡处閹峰煤椤忓秵鏅滈梺鍛婁緱娴滄繐锟???閿熻棄銈稿缁樻媴閸涘﹤鏆堢紓浣割儐閸ㄥ潡寮崘顔芥櫆闁告挆鍜冪闯婵犳鍠楁灙闁糕晜鐗犻幃锟犲即閵忕姷顔愬┑鐑囩秵閸撱劑骞忛敓锟????闂佽法鍠嶇划娆忕暦椤愨挌娲敂閸涱垰�?????闂傚倷绀佹惔婊呭緤娴犲缍栭煫鍥ㄦ礈绾惧吋淇婇婵愬殭妞ゅ孩鎹囧娲川婵犲嫧妲堥梺鎸庢磸閸婃繂顕ｉ幎钘夐唶婵犻潧鍟敓�????婵＄偑鍊栧濠氬Υ鐎ｎ亶鍟呴柕澹懐锛濋悗骞垮劚閹锋垿鐓渚囨闁绘劖褰冮弳锝夋煙椤旂晫鐭掗柟绋匡攻缁旂喖鍩為崹顔碱潎闂佸搫鑻粔鐟扮暦椤愶箑绀嬮柤绋跨仛閺嗕即姊绘担鍛婃儓闁瑰嘲顑嗙粋宥夘敂閸曞灚缍庡┑鐐叉▕娴滄粎绮绘导鏉戠閺夊牆澧介幃濂告煟閿濆娑фい顏勫暣婵℃儼绠涢幘鑸敌掗梻浣规偠閸斿宕￠幎鏂ゆ嫹?閿熻棄鈻庨幒鏃傛澑闂佸湱铏庨崹閬嶅棘閳ь剟姊婚敓锟???濞煎骞忛敓�?????闂佽法鍠撻弲顐ょ不閿燂拷???闂傚倸鍊搁崐鐑芥嚄閸撲礁鍨濇い鏍ㄧ箖閹冲矂鏌ｉ悢鍝ョ煁婵犮垺锕㈠畷顖炲箻椤旇�?鍋撻敓锟???瀵噣宕奸锝嗘珖闂備焦瀵у濠氬疾椤愶箑鍌ㄥù鐘差儐閳锋垿鏌熺粙鍨劉缁惧墽鏁婚弻娑虫�??閿熺瓔鍋呭畷�?勬煥閻曞倹锟?????婵犵妲呴崑鍛崲閸繄鏆︽繛宸簼閸婄兘鏌涘┑鍡楊�?妞ゆ挻妞藉娲箰鎼粹懇鎷荤紓渚囧櫘閸ㄨ泛顕ｉ弻銉ョ厸闁告侗鍠掗幏娲煥閻曞倹锟???????闂傚倷鑳舵灙闁挎洏鍎甸獮鎰板箚瑜夐弸搴ㄦ煏韫囧�????閿熶粙宕戦妸鈺傜厱婵炴垶鈽夐崼銉ョ婵炲樊浜濋埛鎴︽煕濞戞﹫鍔熼柍钘夘樀閺屻劑寮村Ο鍝勫Б婵炲瓨绮岄幉鈽呮嫹?閿燂�??锟藉亹閳ь剚绋掗�?�鍥�?储娴犲鈷戦柛鎰�?级閹牓鏌ㄩ弴姗堟嫹?閿熶粙骞冮敓�????閺佸啴宕掑☉姘妇闂備胶纭堕崜婵喢哄⿰鍩跺洭鏁冮崒娑氬帗闁荤姴娲﹂悡锟犲矗閸曨剦娈介柣鎰彧閼板尅锟???閿熻姤娲�?敃銏ゅ箠閻樿鍨傛繛鎴灻兼竟鏇㈡⒑閸撹尙鍘涢柛鐘冲浮瀵劍绂掞拷?锟筋偆鍘介梺褰掑亰閸樼晫绱為幋锔界厽闊洢鍎抽悾鐢告煛锟??瀣М闁诡喓鍨藉鍫曞箣閻樿京�?勫┑掳鍊楁慨鐑藉磻濞戞碍宕叉俊顖濇閺嗭附銇勯幇鍓佺暠閿燂拷?鐎ｎ喗鏅搁柨鐕傛�?????濠电姷顣槐鏇㈠磻閹达箑纾归柡宓本缍庢繝鐢靛У閼瑰墽澹曟繝姘厵闁硅鍔﹂崵娆撴煕濮橆剛绉洪柡灞界Х椤т線鏌涢幘瀵告噰闁糕晝鍋ら獮�?�晜閽樺鍋撻悜鑺ョ厾缁炬澘宕晶顖炴煕閺囥垻鐣烘慨濠呮缁瑩宕犻埄鍐╂毎缂傚�?�娴囬褔鎮ч崱娑欏仼鐎瑰嫭鍣村ú顏嶆晜闁告洦鍘兼慨锔戒繆閻愵亷�????閿熺晫鏁繝鍥ㄢ挃鐎广儱妫涢々鍙夌節婵犲倻澧涢柣鎾寸懇閹鎮介惂鏄忣潐缁傛帡鏁冮崒娑虫�??閿熻姤鎱ㄥ鍡楀箺閿燂拷?鐎ｎ喗鐓涢敓�????閳ь剟宕伴弽褏鏆︽繛鍡樻尭鍥撮梺绯曞墲椤ㄥ繑�?�奸敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣插亾閿濆應妲堥柕蹇曞Х椤︽澘顪冮妶鍡欏缂佸鍨剁粋鎺撶附閸涘ň鎷哄┑顔炬嚀濞村嫰骞忛敓�?????闂佽法鍠嶇划娆忕暦瑜版帩鏁嗗ù锝勮濞叉悂鎮峰⿰鍛暭閻㈩垱顨婇幃鈥斥枎閹惧鍘介梺鐟邦嚟閸婃牠骞嬮悩杈╁墾闂佹眹鍨归幉锟犳偂閺囥垺鐓涢柛灞剧箖绾爼鏌涢埡�?�М闁哄瞼鍠栭�?�娆戠驳鐎ｎ偆鏆梻浣烘�?瀵爼骞愰幎鑺ユ櫢闁跨噦�??????闂備浇妫勶拷?锟筋剟濡剁粙娆炬綎闁惧繐�?遍惌娆撴煕瑜庨�?�鍛嚕閻楀牏绠鹃悗娑欘焽閻鏌涙惔锝呭付閾荤偤鏌ｉ弬娆炬疇婵炴挸顭烽弻鏇㈠醇濠靛浂妫ゆ繝�???鍥︽喚闁哄本绋撻�?顒婄秵閸嬪棗煤閹绢喗鐓欐い鏇炴閿燂�???闂佽法鍠曡閿燂�??娴犲鍊甸柨婵嗙凹缁ㄨ姤銇勯敓锟???閸旀洟鍩為幋锔斤�??锟介柛銉㈡櫇鏍￠梻浣告啞閹稿鎮烽敂鐣屸攳濠电姴娲﹂崵鍐煃閸濆嫬鏆熼柨娑欑矒濮婅櫣绱掑Ο蹇ｄ邯楠炴牠顢曢敓锟???鐟欙箓鏌涢敂璇插箻缁炬儳銈稿鍫曞醇濞戞ê顬堝┑鐐存儗閸犳濡甸崟顖氼潊闁挎稑瀚崳褔姊猴�??锟界媭鍤欓梺甯秮楠炲啫鈻庨幙鍐╂櫌闂佺ǹ鏈花浠嬪Ψ閳哄�?�鎷绘繛杈剧悼閻℃棃宕靛▎鎾达拷?锟芥繛鎴炲笚濞呭﹪鏌熼搹顐ょ畺闁靛牞缍佸畷锟??濡搁獮顖氭噽绾惧ジ鎮楅敐搴�?�航闁稿簺鍎茬换娑㈠礂閼测晛顫х紓浣虹帛缁嬫垿顢欒箛娑辨晩闁煎鍊曢崵顒勬⒒娴ｈ鍋犻柛濠冪墱閺侇噣鏁撻悩鑼舵憰闂佸搫娲㈤崹褰掓煁閸ャ劎锟??闂傚牊绋掗幖鎰版煛閸涱剛鐭欐慨濠冩そ楠炴劖鎯旈敐鍥╂殼闂備浇顕栭崰鏍ь焽閿熺姴绠栭柣鎴ｆ缁犮儵鏌涢幇顖氱毢濠�?屽灦濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犲ù鐓庣摠閻撴洟鏌熼悜妯诲碍缂佹甯￠弻宥囨嫚閸欏鏀紓浣哄У閻╊垰顕ｉ幘顔藉亜闁告挻褰冮弲顓熺節閻㈤潧啸闁轰焦鎮傞弫鎾绘晸閿燂拷??婵犵數鍋�?崠鐘诲炊閵娿儰缃曢梻浣告啞娓氭宕㈤幖浣歌摕闁挎柨顫曟禍婊堢叓閸ャ劍灏靛褎鐩弻娑虫嫹?閿熺獤鍐ㄢ拤缂備胶绮惄顖氱暦閸楃�?�鐔煎礂閻撳孩鐝紓鍌氾�??锟界粈锟??顢栭崨杈炬嫹?閿熶粙鎮滈挊澶庢憰闂佹寧绻傚Λ娆撳磿閻斿吋鐓忥�??锟界増鐩�?�锕傛惞鎼淬垻锟??婵炲牆鐏濋弸娑㈡煥閺囨ê濡奸柍璇茬Ч閺佹劖寰勬繝鍕瀫闂備礁�?遍搹搴ㄥ窗閺嶎偆鐭嗛悗锝庡亖娴滄粓鏌熸导瀛樻锭濞存粍绻冮妵鍕Ψ閵夘喖鍓伴梺�?�狀潐閸ㄥ潡骞冮埡鍜佹晝闁挎繂鎷嬮埀�???绻樺娲川婵犲啰顦ラ梺璇茬箲锟??鎼佸箖閸ф鏅搁柨鐕傛�??闂佽鍠楅�?�鍛村煝閹捐鍨傛い鏃傛櫕娴滃爼姊绘担铏瑰笡闁圭⒈鍋嗛幑銏犫攽鐎ｎ偄浠掗梺璺ㄥ櫐閿燂�???閻庢鍠曠划娆愪繆閹间焦鏅搁柨鐕傛嫹?濡炪倕�?�╅幑鍥ь潖濞差亝顥堥柍杞拌兌濡诧綁姊洪崨濠庣劷闁告鍥舵晪闁挎繂顦粻锟??鏌ら幁鎺戝姉闁归绮换娑欐綇閸撗呅氬┑鐐叉嫅缁插潡寮灏栨婵炲棙鍨归鏇㈡⒑閸涘﹦鎳冩い锕�?哺閺呭墎鍠婃径�?��??闂佽法鍠曟慨銈吤洪敓�????瀹曟繂顫滈埀顒佷繆閻㈢ǹ绠涢柡澶庢硶椤斿﹪姊虹憴鍕姢闁宦板姂椤㈡棃鎮㈤崗灏栨嫽婵炶揪�???婵倗娑甸崼鏇熺厱闁挎繂绻掗悾鐢告煥閻曞倹锟????????
        .ren(backend_dcache_ren),
        .wen(backend_dcache_wen),
        .writen(backend_dcache_writen),
        .vaddr(backend_dcache_addr),
        .write_data(backend_dcache_write_data),
        .llw_to_dcache(llw_to_dcache),
        .scw_to_dcache(scw_to_dcache),

        //trans_addr to dcache
        .ret_data_paddr(ret_data_paddr),
        .duncache_en(duncache_en),
        .is_exception_execute1_i(is_exception_execute1),

        .data_addr_trans_en(data_addr_trans_en),
        .data_tlb_found(data_tlb_found_out),
        .data_tlb_v(data_tlb_v_out),
        .data_tlb_d(data_tlb_d_out),
        .csr_plv(csr_plv),
        .data_tlb_plv(data_tlb_plv_out),

        .icacop_en(icacop_en),
        .dcacop_en(dcacop_en),
        .cacop_mode(cacop_mode),
        .cache_cacop_vaddr(cache_cacop_vaddr),
        .cache_axi_write_pre_ready(cache_axi_write_pre_ready),

        // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠楅悷鈺侇嚕閸洖鍨傛い鏇炴噹濞堫參姊婚崒姘炬�??閿熶粙宕愰幖浣哥９闁绘垼濮ら崐鍧楁煥閺囩儑锟???閿熺晫绮婚弽顓熺厱妞ゆ劧绲鹃敓锟???缂佺偓鍎冲锟犲蓟閿濆绠ｉ柣鎴濇閸斿嘲顪冮妶鍌涙珔鐎殿喖澧庨幑銏犫攽閸モ晝鐦堥梺绋挎湰缁矂路閳ь剟姊绘担鍛佃顨ラ崫銉х煋鐟滅増甯掗拑鐔兼煥濠靛棭妲哥紒鐙呯秮閺岋綁骞囬敓�????閺嗙偟绱掗鑲┬ょ紒顔碱儏椤撳ジ宕ㄩ鍕闂備礁澹婇崑鍡涘窗閹捐鐭楅柛鈩冪⊕閳锋垿鏌涘┑鍡楊仼闁哄棙鐟︾换娑㈠级閹存績鍋撻崹顔炬殾闂傚牊绋堥弸搴ㄦ煙鐎涙ɑ鐓ュù婊呭亾缁绘盯宕煎┑鍫滆檸濠电偛鎳忛敃銏ゅ蓟濞戙垺鏅查煫鍥ㄦ礈琚﹂柣搴㈩問閸犳牠鈥﹂悜钘夊瀭闁诡垎鍛闂佹悶鍎崝宥夋偩閻戣姤鈷戦悹鍥ㄥ絻閸よ京绱撳鍛棦鐎规洘绮岄埥澶娾攦閹冪�?闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊椤掑鏅梺鍝勭▉閸樿偐绮ｅΔ鍛厵闁绘垶锕╁▓鏃堟煟閵堝洤浜剧紒缁樼箖缁绘繈宕掑顓犱壕闂備胶绮敮濠勫垝濞嗘挻鍋傛い鎰剁畱閻愬﹪鏌曟繛鍖℃�??閿熺晫鎹㈤敓�????濮婄儤娼幍顕呮М闂佸摜鍣ラ崹鑸典繆閻㈢ǹ绀嬫い鏍ㄦ皑閿燂拷?闂備礁鐤囧銊╂嚄閼哥數顩峰┑鍌氭啞閳锋帒鈹戦悩鑼闁伙絽鐏氶幈銊︾節閸屻倗鍚嬮悗瑙勬礃鐢帡锝炲┑�?�垫晞闁芥ê顦竟鏇㈡⒑缂佹ê鐏卞┑顔猴�??锟藉畷鐢稿礋椤栨稓鍘遍梺瑙勫礃鐏忔瑩藝閿曞�?�鐓曢柕濠忓缁犳牠鏌曢崶褍顏�??锟筋喕绮欓�?�鏇綖椤撶姵宕熺紓鍌氾�??锟介懗鑸垫叏閹惰棄锟??闁规儼妫勯拑鐔兼煟閺傚灝鎮戦柍閿嬪浮閹鎮介惂鏄忣潐娣囧﹥绂掞�??锟筋�?鎷虹紓浣割儐椤戞瑩宕曡箛鏂讳簻闁瑰瓨绻嶉敓锟???閻庢鍠栭�?�鐑藉箖閵忋倕绀傜痪顓㈡敱閿燂拷??闂佽法鍠曟慨銈夊Φ閸曨垰绠抽柛鈩冦仦婢规洖鈹戦悩顐ｅ�?�閻忕偟鏅禒鎼佹⒑閸濆嫭婀伴柣鈺婂灡娣囧﹪宕奸弴鐐诧拷?锟藉┑鈽嗗灣閳峰牆危瑜版帗鈷掑ù锝呮啞閹牓鏌￠崼顐㈠⒋闁诡垰瀚伴、娑㈡�?�闂堟稓銈﹂梻浣规偠閸庢椽宕滈敃鍌氭瀬闁搞儺鍓氶悡鐔告叏閿燂�??濡寮稿☉妯忓綊鎮崨顖滄殼濠殿喖锕︾划顖炲箯閸涱垳鐭欐繛鍡欏亾椤ユ垿姊绘担鍛靛綊顢栭崱娆愭殰婵°�?�鍟伴惌澶涙�??閿熷鍎遍ˇ浠嬪极閸岀偞鐓曟い鎰剁悼缁犳岸鏌熼懞銉︾闁宠鍨块幃娆撳级閹寸姳鎴烽梻浣虹�?�閺呮冻�????閿熻姤婢�?锝夘敃閿燂�??�???鍐┿亜閺冨�?�娅曢柛姗嗕邯濮婃椽宕滈幓鎺嶇凹缂備浇顕ч崯鏉戠暦閸愯娲敂閸涱垰骞楅梻濠庡亜濞层�?�霉妞嬪海鐜婚柡鍐ｅ亾闁逛究鍔嶇换婵嬪礃閳瑰じ铏庨柣搴ゎ潐濞插繘宕濆鍥ㄥ床婵炴垯鍨圭粻铏�?闂堟稒鍤囬柛瀣殜濮婅櫣鎷犻垾铏亶闂佹寧纰嶉妵鍕敃閿濆洨鐤勫銈冨灪閿曘垽骞冮埡鍜佹晝闁挎繂妫欏▓鐓庘攽閻樺灚鏆╁┑顔惧厴�?�偊宕ㄦ繝鍐ㄥ伎闂佸搫顦伴崵姘洪鍛珖闂佺ǹ鏈銊╂晬濞嗘劒绻嗛柣鎰▕閸庡繒绱掗妸銉у煟鐎规洘鍨块獮妯肩磼濡桨鐢婚梻浣告惈椤︿即顢栧▎寰稑鐣濋崟顑芥嫼闂佸憡绺块崕杈ㄧ墡闂備胶绮〃鍫熸叏閹绢喗鍋╋拷?锟藉嫭澹嬮崼顏堟煕椤愩�?�鏋庡ù婊堜憾濮婃椽宕滈幓鎺嶇凹缂備緡鍠栧ù椋庡垝鐠囧樊娼╅柤鍝ヮ暯閹锋椽姊婚崒姘卞�?缂佸鎸婚弲鍫曞即閻旇櫣顔曢柣蹇曞仜閸嬪﹪骞忛敓�?????闂佽法鍠嶇划娆撳箖瑜庨幆鏃堝Ω閿旇�?�藉┑鐐舵彧缁插潡鎮洪弮鍫濆惞闁告劦鍠楅悡鏇㈡煟濡櫣锛嶅褏鏁搁埀顒冾潐濞叉﹢宕濆▎鎾跺祦闁哄秲鍔嶆刊鎾煟閻旂⒈鏆掗柟顕嗙秮濮婄粯鎷呴搹鐟扮闂佹悶鍔庨崢褑鐏嬮梺鍛婃处閸ㄧ晫绱為弽顓熺厱婵炴垶顭囬幗鐘绘煟閹惧磭绠婚柡灞剧洴椤㈡洟鏁愰崶鈺冩毇闂備線娼婚敓�????濠殿喓鍊濋弫鎾绘晸閿燂拷????闂佹眹鍩勯崹杈╂暜閿熺姴鐏抽柡鍐ㄧ墕�???鍐┿亜閺傛寧顫嶇憸鏃堝蓟濞戙垹鐒洪柛蹇ラ檮锟??鎼佺嵁韫囨梻�???婵﹩鍘搁幏娲⒑閸涘﹦绠撻悗姘煎幗閸掑﹥绺介崨濠勫幈闁诲函缍嗘禍宄邦啅閵夆晜鐓熼柨婵嗘搐閸樻挳鏌ㄩ悤鍌涘?闂備線娼ч悧鍡涘箠鎼达絿鐜绘繛鎴炵懅閿燂拷?闂佹眹鍨藉褍鐡梺璇插閸戝綊宕抽敐澶涙嫹?閿熻棄鈻庨幘鍐插祮闂�?潧楠忕槐鏇㈠储閸涘﹦�???闁靛骏绲剧涵楣冩煥閺囶亪妾柡鍛埣瀵挳鎮滈崱娆忔暩闁荤喐绮岀换妯侯嚕閺屻儺鏁冮柕鍫濇噹閻忓﹪姊洪崫鍕殭闁绘绮撳顐﹀幢濡炴洖缍婇弫鎰板川椤撶噦锟???閿熺晫绱撴担闈涘妞ゆ泦鍥锋�??閿熶粙宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣鍖栭弴鐔哥彅闁诲孩鍑归崜娆忕暤閸曨垱鈷戠憸鐗堝笚閿涚喖鏌ｉ幒鐐电暤闁诡噯绻濋幃銏ゅ礂閼测晛寮虫繝鐢靛█濞佳兾涘▎鎾抽棷閻熸瑥�?�换鍡涙煙缂佹ê淇柣鎾炽偢閺岋�??锟界暆鐎ｎ剛袦闂佽桨鐒﹂崝娆忕暦閸楃偐鏋庨柟瀵稿У濠㈡牠姊虹拠鍙夊攭妞ゎ偄顦叅婵犲﹤鐗嗙粣妤呮煛瀹ュ骸寮块柟鍑ゆ�??闂佽法鍠曞Λ鍕亙闂佸憡渚楅崢楣冩晬濠婂啠�?芥い�???鏋绘笟娑㈡煕閹惧娲存い銏∩戠缓浠嬪川婵炵偓瀚介梺璺ㄥ櫐閿燂�???????闂傚倷鑳剁划顖滄暜椤忓棛涓嶉柟鎯х－閺嗭箓鏌￠崶銉ョ仼閿燂�??閸愵喗鍋″ù锝囨焿閸忓矂鏌熼搹顐ｅ磳闁挎繄鍋涢埞鎴�?醇閻旈锛忛梻浣瑰劤缁绘帒鈻嶉姀銏☆潟妞ゆ洍鍋撴慨濠呮閹风�?骞撻幒鎴炵槪缂傚倸鍊哥粔鏉懳涘┑鍡欐殾闁瑰墎鐡旈敓锟????闁诲孩顔栭崳�???宕戞繝鍌滄殾闁圭儤顨嗛崐鐑芥倵閻㈢櫥褰掔嵁閸喍绻嗛柣鎰典簻閳ь剚鐗犲畷婵嬫晝閸屾氨锛涢梺鍛婃处閸撴艾鈻嶉悩缁樼厵婵炲牆鐏濋弸銈囩棯閹佸仮闁诡喗顨婇弫鎰償濠靛牊鏅肩紓鍌欒兌婵娊宕￠幎钘夎摕鐎广儱娲﹂崰鍡涙煕閺囥劌浜炲ù鐓庣焸濮婅櫣鎷犻垾铏亐闂佸搫鎳忕换鍕ｉ幇鏉跨闁瑰啿纾崰鎰崲濠靛棭娼╂い鎾跺枑椤斿啫鈹戦悩娈挎殰缂佽鲸娲熷畷鎴﹀箣閿燂拷?绾惧綊鏌″搴�?�箹闁搞劌鍊块弻锝夊閳惰泛�?辩划濠氭偐缂佹鍘甸梻渚囧弿缁犳垿宕拷?锟芥ü绻嗛柟缁樺笧婢э箓鏌�?�畝瀣М濠殿喒锟????闂傚倷鑳剁划顖滄暜閹烘鍊舵慨妯挎硾妗呴梺鍛婃处閸ㄦ壆绮婚幎鑺ョ厵閻庢稒顭囩粻銉ッ归悩鑽ょ暫婵﹥妞介獮搴ㄦ嚍閵夛附娈搁梻浣规偠閸斿苯锕㈤崡鐐嶏綁骞囬弶璺啋闁诲孩绋掗敋妞ゅ孩鎸荤换婵嗏枔閸喗鐏嶉梺绯曟櫅閻�?﹦绮嬪鍛�?閻庯綆浜為悿鍕⒑闂堟单鍫ュ疾濞戙垺鍊峰┑鐘插暔娴滄粓鏌熼崫鍕ラ柛蹇撶焸閺屾稑螣閸︻厾鐓撳┑鈽嗗亜閹虫﹢銆�?弴銏�?潊闁炽儲鍓氬Σ閬嶆⒒娴ｅ憡鎯堥悶姘煎亰瀹曟繈骞嬪┑鍫熸濡炪�?�鍔ч梽鍕磹缂佹ü绻嗘い鏍仦濞呮粎绱掗妸銉吋婵﹥妞藉Λ鍐ㄢ槈濮樿京鏆伴梻浣虹�?�閺呮冻�????閿熸垝鍗抽悰顕嗘�??閿熺瓔鍠楅崑鎰版煕閹邦厼绲荤紒銊ｅ劜缁绘繈鎮介棃娑掓瀰濠电偘鍖犻崗鐐洴椤㈡﹢鎮滈崱娆忓Ш闂備礁鍟块幖顐﹀磹閼哥數顩叉繝濠傜墛閻撴瑩鏌熼鍡楄嫰閿燂拷??闂傚倷娴囬褝锟???閿熻В鏅滅粚閬嶅传閸曞孩鐩畷鐔碱敍濮樺崬骞嬮梻浣侯攰閹活亪姊介崟顖氱９闁绘垼濮ら悡鐘绘煙闂傚鍔嶆繛鎳峰嫮绠鹃柟鍐插槻閹虫劗澹曢挊澹濆綊鏁愰崶銊ユ畬缂備浇灏欑划顖滄崲閿燂拷?????闂備椒绱徊鍧楀礂濡警鍤曢柟缁㈠枛椤懘鏌ｅΟ鑽ゅ灩闁告劕澧介崬鐢告煟閻樼儤顏犻悘蹇嬪妼椤斿繘濡烽埡鍌滃幍濡炪�?�鐗楃划灞剧鏉堛劍鍙忓┑鐘插暞閵囨繈鏌＄仦鑺ュ殗闁诡喗鐟╅幊鐘垫崉娓氼垯绱�?繝鐢靛Л閹峰啴宕橀鍛枛闂備緤锟???閿熺晫鈹掗柛鏂跨Ф閹广垹鈹戯拷?锟筋亞顦ㄩ梺宕囨�?閵囨﹢鎼规惔顫箚闁靛牆娲ゅ暩闂佺ǹ顑囬崑銈夊箖瑜旈幃鈺冩嫚閼碱剛鏆繝鐢靛Т閿曘�?�鎮ч崱娑欙拷?锟藉┑鐘叉处閻撳繐鈹戦悙鑼虎闁告梹鎸抽弫鎾绘晸閿燂�?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殘閳ь剙绠嶉崕鍗灻洪妶澶婂瀭婵犻潧娲ㄧ粻楣冩煕閳╁叐鎴犱焊椤撶姷纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍣ｅ畷鐓庘攽閸垺姣囬梻鍌欑閸熷潡骞栭�???鐤い鏍ワ拷?锟介敓锟????闂佽法鍠曟慨銈呯暆閹间礁钃熸繛鎴炃氶弸搴ㄧ叓閸ラ绋诲Δ鏃堟⒒閿燂�??閳ь剛鍋涢懟顖涙櫠婵犳碍鐓曢柟鎹愭硾閺嬪孩銇勯銏㈢閻撱倖銇勮箛鎾村櫣濞寸媭鍙冨娲传閸曞灚笑缂備降鍔戞禍鍫曠嵁閹版澘�?冩い蹇撴閿涙繃绻涢幘纾嬪婵炲眰鍊曢埢宥咁潨閳ь剟寮诲☉銏犖╅柕濠忓閵嗘劕顪冮妶鍡樼┛缂傚秳绀�?锝嗙節濮橆儵銊╂煏婢诡垰鑻弲锝嗙�?閻㈤潧浠╅柟娲讳簽�?�板﹪鎸婃径娑虫�??閿熶粙姊洪敓�????缁夋挳鎯屽Δ鍛厱闁斥晛鍟伴埊鏇㈡煃闁垮鐏╃紒杈ㄦ尰閹峰懘鎯傞崨濠傤�????闂傚倸鍊烽懗鑸电仚闂佹寧娲忛崐鏇㈡晝閵忋倖鐒硷拷?锟姐儱鎳愰崝�???顪冮妶鍡楃瑐闁煎啿鐖煎畷顖炲蓟閵夛妇�??????
        .rdata(dcache_rdata),
        .rdata_valid(dcache_backend_rdata_valid), 
        .sc_cancel(sc_cancel_to_backend),
        .uncache_out(uncache_out),
        .dcache_is_exception(dcache_is_exception),
        .dcache_exception_cause(dcache_exception_cause),   
        .dcache_ready(dcache_ready),  
        .data_fetch(data_fetch),

    //to write BUS
        .dev_wrdy(dev_wrdy_to_cache),      
        .cpu_wen(dcache_wen),        
        .cpu_waddr(dcache_awaddr),      
        .cpu_wdata(dcache_wdata),      
    //to Read Bus
        .dev_rrdy(dev_rrdy_to_cache),       
        .cpu_ren(dcache_ren),        
        .cpu_raddr(dcache_araddr),      
        .dev_rvalid(dcache_rvalid),     
        .dev_rdata(dcache_axi_data_block),
        .ren_received(dcache_ren_received),
    //duncache to cache_axi
        .uncache_rvalid(duncache_rvalid),
        .uncache_rdata(duncache_rdata),
        .uncache_ren(duncache_ren),
        .uncache_raddr(duncache_raddr),

        .uncache_write_finish(duncache_write_finish),
        .uncache_wen(duncache_wen),
        .uncache_wstrb(duncache_wstrb),
        .uncache_wdata(duncache_wdata),
        .uncache_waddr(duncache_waddr)  
    );
        
    addr_trans u_addr_trans
    (
        .clk(aclk),
        .asid(asid_in),
        //inst addr trans   鎸囦护鍦板潃杞�?
        .inst_fetch(inst_rreq),
        .inst_vaddr(inst_addr1),
        .inst_vaddr_plus(inst_addr2),

        .not_same_page(not_same_page),
        .inst_uncache_en(iuncache_en),
        .inst_paddr_out(inst_paddr),
        
        .inst_tlb_found_out(inst_tlb_found),
        .inst_tlb_v_out(inst_tlb_v),
        .inst_tlb_d_out(inst_tlb_d),
        .inst_tlb_mat_out(inst_tlb_mat),
        .inst_tlb_plv_out(inst_tlb_plv),
        .inst_addr_trans_en_out(inst_addr_trans_en),
       
        //data addr trans   鏁版嵁鍦板潃杞�?
        .data_fetch(data_fetch | is_tlbsrch),
        .data_vaddr(backend_dcache_addr),
        .dcacop_en(dcacop_en),
        .cacop_mode(cacop_mode),

        .data_uncache_en(duncache_en),
        .data_paddr_out(ret_data_paddr),

        .tlbfill_en(tlbfill),
        .tlbwr_en(tlbwr),

        .data_tlb_found_out(data_tlb_found_out),
        .data_tlb_index_out(data_tlb_index_out),
        .data_tlb_v_out(data_tlb_v_out),
        .data_tlb_d_out(data_tlb_d_out),
        .data_tlb_mat_out(data_tlb_mat_out),
        .data_tlb_plv_out(data_tlb_plv_out),
        .data_addr_trans_en_out(data_addr_trans_en),
 
        //tlbwi tlbwr tlb write
        .rand_index(rand_index),
        .tlbehi_in(tlbehi_in),
        .tlbelo0_in(tlbelo0_in),
        .tlbelo1_in(tlbelo1_in),
        .tlbidx_in(tlbidx_in),
        .ecode_in(ecode_in),


        //tlbr tlb read
        .tlbehi_out(tlbehi_out),
        .tlbelo0_out(tlbelo0_out),
        .tlbelo1_out(tlbelo1_out),
        .tlbidx_out(tlbidx_out),
        .asid_out(asid_out),

        //invtlb 
        .invtlb_en(invtlb),
        .invtlb_asid(invtlb_asid),
        .invtlb_vpn(invtlb_vpn),
        .invtlb_op(invtlb_op),
        //from csr

        .csr_plv(csr_plv),
        .csr_dmw0(csr_dmw0),
        .csr_dmw1(csr_dmw1),
        .csr_da(csr_da),
        .csr_pg(csr_pg),
        .csr_datm(csr_datm),
        .csr_datf(csr_datf)
    );

    axi_interface u_axi_interface(
        .clk(aclk),
        .rst(rst),
    //connected to cache_axi
        .cache_ce(axi_ce_o),
        .cache_wen(axi_wen),   
        .cache_wsel(axi_wsel),      
        .cache_ren(axi_ren),         
        .cache_raddr(axi_raddr),
        .cache_waddr(axi_waddr),
        .cache_wdata(axi_wdata),
        .cache_rready(axi_rready),    
        .cache_wvalid(axi_wvalid),     
        .cache_wlast(axi_wlast),      
        .wdata_resp_o(axi_wdata_resp),    
    
        .cache_brust_type(cache_brust_type),  
        .cache_brust_size(cache_brust_size),
        .cacher_burst_length(axi_rlen),
        .cachew_burst_length(axi_wlen),

        .arid(arid),       
        .araddr(araddr),      
        .arlen(arlen),      
        .arsize(arsize),
        .arburst(arburst),
        .arlock(arlock),   
        .arcache(arcache),   
        .arprot(arprot),   
        .arvalid(arvalid),       
        .arready(arready),         
    //R闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归崷顓犱笉閻犲洩顥嗚ぐ鎺撴櫜闁割偒鍋呯紞鍫ユ⒑闂堟稒澶勭紒璇插暣婵＄敻宕熼姘兼綂闂佹枼鏅涢崰姘涢崘顔斤�??锟介悷娆忓绾炬悂鏌涢敓�????閸ㄥ潡濡存担鑲濈喓鎮伴埄鍐╂澑闂備礁澹婇崑鍡涘窗閹邦儷鎺撴償閵婏腹鎷婚梺绋挎湰閻旑剟骞忛敓锟????闂佽法鍠嶇划娆忕暦閹邦収妲归幖杈剧悼閿燂�????婵°�?�濮烽崑鐐烘偋閻樹紮�????閿熶粙寮村杈┬㈤梻浣规偠閸庢椽宕滃▎鎴犱笉闁靛�?璐熸禍婊堟煛閸愵煉锟???閿熶粙宕甸埀顒佺箾鐎涙鐭婂褏鏅Σ鎰板箳閹宠櫕姊归幏鍛偘閳╁喚娼斿┑鐘垫暩閸嬬偛顭囧▎鎾崇９闁割煈鍣�?崵鏇熴亜閹板墎鎮肩紒�???鍋撻梻浣规偠閸庮垶宕濇惔銊ュ偍闁瑰墽绮崑鈩冪節婵犲倸顏柣顓熷笧閳ь剝顫夊ú妯煎垝閹捐绠栭柕蹇ョ磿闂勫嫬顭跨捄渚剳缂佸鑳剁槐鎾诲磼濮橆兘鍋撻悜鑺ワ拷?锟介柨鏇氱劍閹冲苯鈹戦悩鎰佸晱闁搞劑浜堕獮鎰板箮閽樺鎽曢梺闈涚墕椤︻垳绮婚幒妤佺厵闁绘垶锚閻忋儱鈹戦鍝勭伈婵﹥妞藉Λ鍐ㄢ槈濞嗘ɑ顥ｉ梻浣瑰濞诧附绂嶅⿰鍫稏闊洦鎷嬪ú顏嶆晜闁告粈鐒﹂ˉ鍫ユ⒒娴ｇǹ鏆遍柟纰卞亰瀹曨垶骞忕仦瑙ｅ亾鐎靛摜纾介柛灞捐壘閳ь剛鍏橀幊妤呮嚋閸偄寮块梺姹囧灮鏋紒鐘崇�?閺屾盯濡烽鐓庮潽闂佺ǹ顑嗚摫闁靛洤�?�板锟??宕堕妸褝�???????婵犵數濮烽弫鎼佸磻閻愬搫鍨傞柛顐ｆ礃閸嬶繝鏌ㄩ悤鍌涘�??闂佸疇顕х粔瑙勬叏閳ь剟鏌曢崼婵囶棏闁归攱妞介弻锝夋偐閸忓懓鍩呴梺鍛婃煥閼活垶鍩㈠澶婄�?闁绘鐗忛崢鐢告⒑閸涘﹤鐏熼柛濠冪墵閺佹捇鏁撻敓�???????
        .rid(rid),
        .rdata(rdata),   
        .rresp(rresp),    
        .rlast(rlast),           
        .rvalid(rvalid),       
        .rready(rready),
        .rdata_o(axi_rdata),
        .rdata_valid_o(axi_rdata_valid),         
    //AW闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁诡垎鍐ｆ寖闂佺娅曢幑鍥灳閿燂拷?????婵＄偑鍊曠换鎰板箠韫囨挾鏆﹂柟鎯板Г閳锋垶绻涢懠棰濆殭妤犵偞鐗楁穱濠囶敃閿濆洨鐤勯悗娈垮枛椤攱淇婇幖浣哥厸闁稿本鐭花浠嬫⒒娴ｅ懙褰掑嫉椤掑倻鐭欓柟杈惧瘜閿燂拷???婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙稑鈹戦悙鏉戠亶闁瑰磭鍋ゅ畷鍫曨敆娴ｉ晲缂撶紓鍌欑椤戝棴�????閿熺獤鍥拷?锟芥い鎺戝閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁悗瑙勬礃閸ㄥ潡鐛崶顒佸亱闁割偁鍨归獮妯肩磽娴ｅ搫浜炬繝銏∶悾鐑筋敆娴ｈ鐝风紓鍌欑劍鐪夌紒璇叉閺屻�?�鍠婇崡鐐差潻闂佸憡锚閻°劑骞堥妸锔剧瘈闁告洦鍘肩粭锟犳⒑閻熸澘妲婚柟铏悾鐑藉Ω閿斿墽鐦堥梺鍛婂姂閸斿本绔熷鍥╃＝闁稿本鑹鹃埀顒勵棑缁牊绗熼�?顒勶�??锟介弽顓炵妞ゆ挾鍣ラ崑銊モ攽椤�?枻渚涢柛鎾寸洴�?�娊鏁冮崒娑氬帾闂婎偄娲㈤崕宕囧閹稿簺浜滈柍鍝勫暙閸樻挳鏌熼绛嬫疁闁轰焦鍔栭幆鏂库攽閸喐娅﹂梻鍌欑劍鐎笛呯矙閹烘鍎庢い鏍ㄥ嚬濞兼牠鏌ц箛姘兼綈鐎规洖顦甸弻鏇熺箾閸喖濮曢梺璇茬箣閻掞妇鎹㈠┑鍡忔灁闁割煈鍠楅悘鎾绘⒑鏉炴壆顦︽い顓犲厴閻涱噣宕�?鑺ユ闂佺粯枪鐏忔瑩藝閵娿儺娓婚柕鍫濇閳锋帡鏌￠崪浣镐喊鐎规洏鍨藉畷锟犳倷閳哄�?�鏉搁梻浣虹帛椤洨鍒掗姘ｆ鐟滃孩绌辨繝鍥舵晝闁挎繂瀛╅悿浣割渻閵堝啫鐏俊顐㈠暣閵嗕線寮崼婵嬪敹闂佺粯鏌ㄩ幖顐︾嵁閸儲鈷掑ù锝囨�?椤曟粎绱掔拠璇ф嫹?閿熶粙鐛繝鍥х疀妞ゆ柨澧介悡瀣攽閻愬弶鈻曞ù婊勭箞閺佹捇鏁撻敓锟??????闂佽鍑界紞鍡涘礈濞戙垺鏅柣鏂垮悑閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曞礈瑜忕壕濂告煕濞嗗浚妲归柕鍥ㄧ箘閳ь剚顔栭崰妤勩亹閸愵喖鐓橀柟杈剧畱闁卞洭鏌曡箛瀣仼缂佺姷鏁诲缁樻媴閸涘﹥鍎撻梺鍝ュ櫏閸嬪﹪骞冭缁绘繈宕堕妸銉ょ暗婵犵數鍋為崹鍫曞春閸愵喖纾婚柟鎹愵嚙�???鍌氼熆鐠虹尨姊楀瑙勬礋濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犻弶鍫㈠亾閿燂拷??闂佽法鍠曟慨銈吤洪幋�???�???闁告劕妯婇崵鏇灻归悩宸剾闁轰礁娲弻锝呂熼崹顔炬闂侀潧鐗炵粻鎾愁潖缂佹ɑ濯村�?�姘煎灡閺侇垶姊虹憴鍕仧濞存粎鍋熼崚鎺撶節濮橆剛顓洪梺缁樏敓�????缂佹顦埞鎴︽倷閺夋垹浠ч梺鎼炲妽濡炰粙宕哄☉銏犵婵°�?�鑳堕崢鍗烆渻閵堝棗濮傞柛濠冩礋瀵悂寮�?崼鐔哄帗濡炪倖鐗楃粙鎺旂矆閸愵喗鐓忛柛銉戝喚浼冮悗娈垮櫘閸撶喎鐣疯ぐ鎺濇晪闁告侗鍓涘Λ顖滅磽閸屾熬�????閿熶粙鎳楅崜浣稿灊妞ゆ牗绮嶅畷鏌ユ煕閺囥劌鐏犵紒鎰殔閳规垿鎮╅煫顓℃姉闂佺粯妫�?鏍惞閸︻厾锛滃┑鈽嗗灥閸嬫劖鏅ラ梻鍌氾拷?锟介崐鎼佸磹閻戣姤鏅搁柨鐕傛�???濠碉紕鍋戦崐鏍垂閻㈢ǹ绠犳慨妞诲亾闁绘侗鍠楃换婵嬪磼閵堝棗缂撻梻渚婃�??閿熻棄鑻晶顔姐亜閺囶亞绉い銏℃礋閺佹捇鏁撻敓�?????缂備讲鍋撻柛鎰ㄦ杺娴滄粓鏌￠崘顭掓嫹?閿熶粙骞忛埄鍐闁绘挸鍑介煬顒佹叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚倷鑳堕�?�濠傗枍閺囥垹绠查柛銉墰�?�撲焦淇婇妶鍛櫣闁告濞婇弻鏇＄疀婵犲喛锟???閿熶粙鏌熼柨瀣仢婵﹥妞藉畷銊︾節閸曨厾鏆ら梺璇插閸戝綊宕ｉ崘銊ф殾闁圭儤顨呮儫闂佸啿鎼崐濠氬储闁秵鈷戦梻鍫熻儐瑜版帒纾匡�??锟芥洖娲ㄩ惌鎾寸箾�?�割喕绨奸柣鎾寸洴閹﹢鎮欓悽鍨啒闂佺ǹ瀛╁Λ鎴﹀箯閿燂拷??闂佽法鍠曟慨銈吤洪弽顓熷亯闁稿繘妫跨换鍡樻叏濠靛棛鐒炬俊鏌ョ畺濮婄儤瀵煎▎鎴犳殸闂佺粯顨嗛幐鎼侊綖韫囨梻�???婵﹩鍓涢敍婊冣攽椤旂煫顏勭暦椤掑嫭鏅搁柨鐕傛嫹?缂傚倸鍊搁崐椋庣矆閿燂拷?椤㈡牠宕卞▎鎰闂佺粯鍔欏褔宕瑰┑鍡忔斀闁绘ê寮堕幖鎰版煟閹惧娲撮柡灞剧〒娴狅箓宕滆閸ｎ喚绱撴担鍝勑ｉ柤褰掔畺閳ユ棃宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣绮欓崠鈩冩暰濠电偛寮堕…鍥╁垝鐎ｎ喖绠抽柟瀛樻煥閻楁岸姊洪崨濠冪５闁哄懏鐟ч懞杈╂嫚瀹割喗�?�岄梺闈涚墕閹虫劗绮绘导瀛橈�??锟芥慨妯煎帶婢ц揪�????閿熺瓔鍠楁繛濠囧极閹版澘宸濇い蹇撴噺閺夋悂姊绘担鍝勪缓闁稿氦浜竟鏇㈩敇閵忕姵锟??????闂備礁鎼ú锕傛晪婵犳鍠栭崐褰掑Φ閸曨垰顫呴柨娑樺閿燂拷??闂備胶顢婇崑鎰偘閵夆晛�?堟繝闈涱儏濮瑰弶銇勮箛鎾跺闁抽攱甯￠弫鎾绘晸閿燂拷??????闂傚倷鑳堕崢褔宕幐搴㈡珷閹兼番鍔岀粈鍡涙煙閻戞﹩娈㈤柡浣哥Ч閺岋綁骞囬鐔虹▏婵炲瓨绮撴禍璺侯潖濞差亜浼犻柛鏇ㄥ墮閸嬪秹姊洪幖鐐插闁硅櫕鎸哥叅閻犳亽鍔庣壕浠嬫煕鐏炲墽鎳呮い锔奸檮閵囧嫰骞嬪┑鍥舵＆濡炪�?�鍨洪悧鏇㈠煝鎼淬劌绠婚柛鎰�?级閸庮亪姊绘担鍛婃儓婵炲眰鍨藉畷鐟懊洪鍕紱闂佹寧绻傞ˇ浼存偂閺囥垺鐓忓鑸电�?�閸掓澘鈹戦垾铏仴闁哄本娲熷畷鐓庘攽閸喐鍠栧┑鐑囩到濞层倝鏁冮鍫㈠祦闁规崘顕х粻鎶芥煛閸屾侗鍎ラ柡澶婃憸缁辨捇宕掑▎鎺戝帯缂備緡鍣崹鎶藉箲閵忋倕绀冩い蹇撴噹鎼村﹤鈹戦悩缁樻锭妞ゆ垵鎳愭竟鏇㈠礂閸忕厧寮垮┑鈽嗗灣閸樠呮暜鐠鸿�?�?介柨娑樺閸樺瓨鎱ㄦ繝鍐┿仢鐎规洦鍋婃俊鐑藉Ψ閿旈敮鍋撴ィ鍐┾拺閻犲浄�????閿熻姤鐏堥梺绋匡攻閹�?�鏁愰悙鍓佺杸闁哄啫鍊婚惁鍫濃攽椤旀枻渚涢柛鎾寸洴閺佸秴饪伴崘锝嗘杸闂佺粯鍔曞鍫曀夐悙鐑樼厱闁哄啠鍋撴い銊ワ攻娣囧﹪宕奸弴鐐甸獓闁圭厧鐡ㄩ幐濠氬棘閳ь剟姊绘担铏瑰笡闁告梹娲栬灒濠电姴浼ｉ敐鍥ㄥ枂闁告洦鍘鹃鏇㈡⒑閼测斁鎷￠柛鎾寸懇�?�憡鎯旈妸锔惧幗闂佹寧绻傚ú銈夊储鐎涙﹩娈介柣鎰叀閸欏嫰鏌熷畷鍥т槐濠碉紕鍏�?弫鍌炴偩鐏炵晫鎮奸梻鍌氾�??锟介崐鐑芥嚄閼哥數浠氶梻浣告惈閻楁粓宕滃▎鎿勭稏婵犻潧顑呮儫闂佸啿鎼敃銉╁疾閳哄懏鈷戠紒顖涙礀婢ц尙绱掞�??锟筋偄娴�?柛鈺傜洴楠炲鏁傞挊澶夊寲闂備浇顕栭崢鐣屾暜閹烘挷绻嗛柛蹇氬亹缁犻箖鏌涘☉鍗炴灈濠殿喖绉归弻鈥崇暆閳ь剟宕伴弽褏鏆︽繛鍡樻尭锟??????
        .awid(awid),     
        .awaddr(awaddr),  
        .awlen(awlen),    
        .awsize(awsize),   
        .awburst(awburst),
        .awlock(awlock),   
        .awcache(awcache),
        .awprot(awprot),   
        .awvalid(awvalid),        
        .awready(awready),        
    //W闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁诡垎鍐ｆ寖闂佺娅曢幑鍥灳閿燂拷?????婵＄偑鍊曠换鎰板箠韫囨挾鏆﹂柟鎯板Г閳锋垶绻涢懠棰濆殭妤犵偞鐗楁穱濠囶敃閿濆洨鐤勯悗娈垮枛椤攱淇婇幖浣哥厸闁稿本鐭花浠嬫⒒娴ｅ懙褰掑嫉椤掑倻鐭欓柟杈惧瘜閿燂拷???婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙稑鈹戦悙鏉戠亶闁瑰磭鍋ゅ畷鍫曨敆娴ｉ晲缂撶紓鍌欑椤戝棴�????閿熺獤鍥拷?锟芥い鎺戝閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁悗瑙勬礃閸ㄥ潡鐛崶顒佸亱闁割偁鍨归獮妯肩磽娴ｅ搫浜炬繝銏∶悾鐑筋敆娴ｈ鐝风紓鍌欑劍鐪夌紒璇叉閺屻�?�鍠婇崡鐐差潻闂佸憡锚閻°劑骞堥妸锔剧瘈闁告洦鍘肩粭锟犳⒑閻熸澘妲婚柟铏悾鐑藉Ω閿斿墽鐦堥梺鍛婂姂閸斿本绔熷鍥╃＝闁稿本鑹鹃埀顒勵棑缁牊绗熼�?顒勶�??锟介弽顓炵妞ゆ挾鍣ラ崑銊モ攽椤�?枻渚涢柛鎾寸洴�?�娊鏁冮崒娑氬帾闂婎偄娲㈤崕宕囧閹稿簺浜滈柍鍝勫暙閸樻挳鏌熼绛嬫疁闁轰焦鍔栭幆鏂库攽閸喐娅﹂梻鍌欑劍鐎笛呯矙閹烘鍎庢い鏍ㄥ嚬濞兼牠鏌ц箛姘兼綈鐎规洖顦甸弻鏇熺箾閸喖濮曢梺璇茬箣閻掞妇鎹㈠┑鍡忔灁闁割煈鍠楅悘鎾绘⒑鏉炴壆顦︽い顓犲厴閻涱噣宕�?鑺ユ闂佺粯枪鐏忔瑩藝閵娿儺娓婚柕鍫濇閳锋帡鏌￠崪浣镐喊鐎规洏鍨藉畷锟犳倷閳哄�?�鏉搁梻浣虹帛椤洨鍒掗姘ｆ鐟滃孩绌辨繝鍥舵晝闁挎繂瀛╅悿浣割渻閵堝啫鐏俊顐㈠暣閵嗕線寮崼婵嬪敹闂佺粯鏌ㄩ幖顐︾嵁閸儲鈷掑ù锝囨�?椤曟粎绱掔拠璇ф嫹?閿熶粙鐛繝鍥х疀妞ゆ柨澧介悡瀣攽閻愬弶鈻曞ù婊勭箞閺佹捇鏁撻敓锟??????闂佽鍑界紞鍡涘礈濞戙垺鏅柣鏂垮悑閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曞礈瑜忕壕濂告煕濞嗗浚妲归柕鍥ㄧ箘閳ь剚顔栭崰妤勩亹閸愵喖鐓橀柟杈剧畱闁卞洭鏌曡箛瀣仼缂佺姷鏁诲缁樻媴閸涘﹥鍎撻梺鍝ュ櫏閸嬪﹪骞冭缁绘繈宕堕妸銉ょ暗婵犵數鍋為崹鍫曞春閸愵喖纾婚柟鎹愵嚙�???鍌氼熆鐠虹尨姊楀瑙勬礋濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犻弶鍫㈠亾閿燂拷??闂佽法鍠曟慨銈吤洪幋�???�???闁告劕妯婇崵鏇灻归悩宸剾闁轰礁娲弻锝呂熼崹顔炬闂侀潧鐗炵粻鎾愁潖缂佹ɑ濯村�?�姘煎灡閺侇垶姊虹憴鍕仧濞存粎鍋熼崚鎺撶節濮橆剛顓洪梺缁樏敓�????缂佹顦埞鎴︽倷閺夋垹浠ч梺鎼炲妽濡炰粙宕哄☉銏犵婵°�?�鑳堕崢鍗烆渻閵堝棗濮傞柛濠冩礋瀵悂寮�?崼鐔哄帗濡炪倖鐗楃粙鎺旂矆閸愵喗鐓忛柛銉戝喚浼冮悗娈垮櫘閸撶喎鐣疯ぐ鎺濇晪闁告侗鍓涘Λ顖滅磽閸屾熬�????閿熶粙鎳楅崜浣稿灊妞ゆ牗绮嶅畷鏌ユ煕閺囥劌鐏犵紒鎰殔閳规垿鎮╅煫顓℃姉闂佺粯妫�?鏍惞閸︻厾锛滃┑鈽嗗灥閸嬫劖鏅ラ梻鍌氾拷?锟介崐鎼佸磹閻戣姤鏅搁柨鐕傛�???濠碉紕鍋戦崐鏍垂閻㈢ǹ绠犳慨妞诲亾闁绘侗鍠楃换婵嬪磼閵堝棗缂撻梻渚婃�??閿熻棄鑻晶顔姐亜閺囶亞绉い銏℃礋閺佹捇鏁撻敓�?????缂備讲鍋撻柛鎰ㄦ杺娴滄粓鏌￠崘顭掓嫹?閿熶粙骞忛埄鍐闁绘挸鍑介煬顒佹叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚倷鑳堕�?�濠傗枍閺囥垹绠查柛銉墰�?�撲焦淇婇妶鍛櫣闁告濞婇弻鏇＄疀婵犲喛锟???閿熶粙鏌熼柨瀣仢婵﹥妞藉畷銊︾節閸曨厾鏆ら梺璇插閸戝綊宕ｉ崘銊ф殾闁圭儤顨呮儫闂佸啿鎼崐濠氬储闁秵鈷戦梻鍫熻儐瑜版帒纾匡�??锟芥洖娲ㄩ惌鎾寸箾�?�割喕绨奸柣鎾寸洴閹﹢鎮欓悽鍨啒闂佺ǹ瀛╁Λ鎴﹀箯閿燂拷??闂佽法鍠曟慨銈吤洪弽顓熷亯闁稿繘妫跨换鍡樻叏濠靛棛鐒炬俊鏌ョ畺濮婄儤瀵煎▎鎴犳殸闂佺粯顨嗛幐鎼侊綖韫囨梻�???婵﹩鍓涢敍婊冣攽椤旂煫顏勭暦椤掑嫭鏅搁柨鐕傛嫹?缂傚倸鍊搁崐椋庣矆閿燂拷?椤㈡牠宕卞▎鎰闂佺粯鍔欏褔宕瑰┑鍡忔斀闁绘ê寮堕幖鎰版煟閹惧娲撮柡灞剧〒娴狅箓宕滆閸ｎ喚绱撴担鍝勑ｉ柤褰掔畺閳ユ棃宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣绮欓崠鈩冩暰濠电偛寮堕…鍥╁垝鐎ｎ喖绠抽柟瀛樻煥閻楁岸姊洪崨濠冪５闁哄懏鐟ч懞杈╂嫚瀹割喗�?�岄梺闈涚墕閹虫劗绮绘导瀛橈�??锟芥慨妯煎帶婢ц揪�????閿熺瓔鍠楁繛濠囧极閹版澘宸濇い蹇撴噺閺夋悂姊绘担鍝勪缓闁稿氦浜竟鏇㈩敇閵忕姵锟??????闂備礁鎼ú锕傛晪婵犳鍠栭崐褰掑Φ閸曨垰顫呴柨娑樺閿燂拷??闂備胶顢婇崑鎰偘閵夆晛�?堟繝闈涱儏濮瑰弶銇勮箛鎾跺闁抽攱甯￠弫鎾绘晸閿燂拷??????闂傚倷鑳堕崢褔宕幐搴㈡珷閹兼番鍔岀粈鍡涙煙閻戞﹩娈㈤柡浣哥Ч閺岋綁骞囬鐔虹▏婵炲瓨绮屽畷顒勫煘閹达附鍋愰悹鍥囧啩绱ｉ梻浣虹帛椤ㄥ懎螞濠靛棛鏆﹂柟鐑橆殔鎯熼悷婊冮叄瀹曚即骞囬悧鍫㈠幐闂佸憡鍔戦崝搴㈡櫠濞戙垺鐓涢柛娑卞枤閿燂拷?闂佸搫鐭夌紞�???鐛崶顒佹櫢闁跨噦锟???濡炪倧绲炬繛濠囧蓟閿濆围闁稿本鐭竟鏇熺節閻㈤潧啸闁轰焦鎮傚畷鎴︽倷閸濆嫬鐎梺鍓插亝濞叉﹢宕戦敓鐘崇叆闁哄洨鍋涢�?�???鎽滄竟鏇㈠箰鎼存稐绨婚棅顐㈡处閹哥偓鏅跺☉銏＄厽闁规崘娉涢弸娑㈡煛锟??瀣М鐎殿噮鍓熼獮鎰償閵忕姵鐎鹃梻鍌欒兌閹虫捇宕崸�???鐤柟缁㈠枛缁犳牠鏌ㄩ悤鍌涘�??濡炪値鍋呯换鍫ュ箖閳╁啯鍎熼柍钘夋妤犲嫭绻濋悽闈浶為柛銊ャ偢閿濈偞寰勬繛鎺撴そ閹垻娑甸柨瀣�??闂佽法鍠曞Λ鍕煡婢舵劕顫呴柍钘夋噺閿燂拷??闂佽法鍠撻弲顐ゆ閹烘鏁婃繛鍡欏亾缂嶅牓鏌ｆ惔銏ｅ闁靛牏枪椤繑绻濆顒傦紲闂佽法鍣﹂敓�??????闂佸綊妫块悞锕傚磻鐎ｎ亖�?介柣妯哄级婢跺嫰鏌涢妶鍛伃闁哄本鐩崺鍕礃閵婏附鍎у┑鐐茬摠缁瞼绱炴繝鍥ц摕闁绘柨鍚嬮崐缁樹繆椤栨繃顏犲ù鐘层偢濮婃椽骞愭惔锝忔�??閿熶粙鏌涢悩宕囧ⅹ妞ゎ偄绻愮叅妞ゅ繐瀚槐鍫曟⒑閸涘﹥澶勯柛锝庡枛椤洭宕奸弴鐔叉嫼缂備礁顑呴悘婵嬵敆閵忋�?�鐓熼柟鍨閿燂拷??闂佽法鍠撻弲顐﹀汲閿曞�?�鐓欓柟娈垮枛椤ｅ吋銇勯妷銉у�?缂佺粯绋撴竟鏇�??閿熺瓔鍋嗚ぐ褍鈹戦埥鍡椾簻闁哥喐娼欓锝夘敃閿燂�??缁犳盯鏌℃径濠勪虎缂佹劖绋戦—鍐Χ閸℃ê鏆楅梺鍝ュУ閸旀瑩銆佸▎鎰窞闁归偊鍘搁幏缁樼箾鏉堝墽鎮奸柟铏崌閺佹捇鏁撻敓锟??????闂傚倷绶￠崜娆戠矓閹绢喖鍨傞柛锟??鍋為悡鏇犳喐鎼搭煉锟???閿熶粙宕拷?锟芥ê鐝旈梺缁樻煥閹芥粎绮绘ィ鍐╃厵閻庣數枪閳ь剚鍨甸～婵堟崉閾忕懓鎽嬪┑鐐差嚟婵挳顢栭崱娑欏亗闁哄洢鍨洪悡鍐煃鏉炴壆顦﹂柡瀣�??锟界换娑㈠醇濞戞浠奸梻鍥ь樀閺岋綁骞�?搹顐ｅ闯闂佺粯甯掗幉锟犲箞閵婏妇�???闁告侗鍣禒鈺冪磽娓氬洤鏋熼柣鐔叉櫅閻ｉ绮欑拠鐐⒐缁绘盯骞嗚婢规洖鈹戞幊閸婃洟宕幍顔碱棜闁兼祴鏅濈壕钘壝归敐鍜佹綘妞ゅ繐鐗婇崐鍫曟煛婢跺鐏嶉敓�????娴犲鐓ユ繛鎴灻顏堟煛閸�?晛澧鹃柟鍑ゆ�??闂佽法鍠曟慨銈吤哄⿰鍫濈獥闁哄稁鍘归�?顑跨閳藉�???閳╁啯鐝抽梻浣虹《閸撴繆鎽梺缁樼箖缁诲牆顫忔繝姘＜婵炲棙甯掗崢锛勭磽娓氬洤娅�?柛銊ф暬楠炴顢曢敂钘変画濠电姴锕わ拷?锟筋厾娆㈤弻銉︾厱闁绘柨鎲＄亸锕傛煙椤旇宓嗘い銏＄懇閺屻劑顢涘顐㈩棜闂備焦�?�х换鍌涱殽閹间礁鍑犻柣鏂垮悑閻撳啴姊洪崹顕呭剰闁诲繆鏅濈槐鎺撴綇閵婏箑闉嶉梺鐟板槻閹冲繘骞堥妸鈺佺闁挎繂鎳嶅Ч锟??鈹戦悙鍙夘棑闁搞劋绮欏濠氬幢濡ゅ﹤鎮戦梺绯曞墲閻熴儵鐛�?崼銉︹拻濞达�?娅ｇ敮娑㈡煥濮樿京妫紓浣靛灩�?�喖鈹戦埄鍐╁唉妤犵偞甯�?��???宕掑⿰鎰簥濠碉紕鍋戦崐鏍ь潖瑜版帩鏁勬繛鍡樻尭閸氳绻涢崱妯诲鞍闁绘挸鍟撮弻�???螣娓氼垱鈻撳┑鈥冲级閹倿骞楅崼鏇熸櫜濠㈣泛顑傞幏娲⒑閸撹尙鍘涢柛锝庡櫍�?�曟洖鈽夊▎鎴狀啎闂佺ǹ绻愰崥瀣煕閹邦喚纾肩紓浣诡焽缁犵偤鏌熼鑽ょ煓婵☆偄鍟埥澶娢旈崘鈺佺婵犵數濮烽�?�钘壩ｉ崨鏉戠；闁告稑鐡ㄩ崑锟犳煃鏉炴媽鍏岄柡鍡檮缁绘繈妫冨☉鍗炲壈闂佽法鍣﹂敓锟????濠碉紕鍋戦崐鏍箰妤ｅ啫绐楅柟閭�?厴閺嬪秹鏌曡箛�?�舵�??閿熶粙鍩涢幋锔藉仯闁诡厽甯掓俊鍏肩箾閸涱喖濮嶉柡�?嬫嫹????
        .wid(wid),     
        .wdata(wdata),  
        .wstrb(wstrb),    
        .wlast(wlast),          
        .wvalid(wvalid),       
        .wready(wready),         
    //闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁诡垎鍐ｆ寖闂佺娅曢幑鍥灳閿燂拷?????婵＄偑鍊曠换鎰板箠韫囨挾鏆﹂柟鎯板Г閳锋垶绻涢懠棰濆殭妤犵偞鐗楁穱濠囶敃閿濆洨鐤勯悗娈垮枛椤攱淇婇幖浣哥厸闁稿本鐭花浠嬫⒒娴ｅ懙褰掑嫉椤掑倻鐭欓柟杈惧瘜閿燂拷???婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙稑鈹戦悙鏉戠亶闁瑰磭鍋ゅ畷鍫曨敆娴ｉ晲缂撶紓鍌欑椤戝棴�????閿熺獤鍥拷?锟芥い鎺戝閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁悗瑙勬礃閸ㄥ潡鐛崶顒佸亱闁割偁鍨归獮妯肩磽娴ｅ搫浜炬繝銏∶悾鐑筋敆娴ｈ鐝风紓鍌欑劍鐪夌紒璇叉閺屻�?�鍠婇崡鐐差潻闂佸憡锚閻°劑骞堥妸锔剧瘈闁告洦鍘肩粭锟犳⒑閻熸澘妲婚柟铏悾鐑藉Ω閿斿墽鐦堥梺鍛婂姂閸斿本绔熷鍥╃＝闁稿本鑹鹃埀顒勵棑缁牊绗熼�?顒勶�??锟介弽顓炵妞ゆ挾鍣ラ崑銊モ攽椤�?枻渚涢柛鎾寸洴�?�娊鏁冮崒娑氬帾闂婎偄娲㈤崕宕囧閹稿簺浜滈柍鍝勫暙閸樻挳鏌熼绛嬫疁闁轰焦鍔栭幆鏂库攽閸喐娅﹂梻鍌欑劍鐎笛呯矙閹烘鍎庢い鏍ㄥ嚬濞兼牠鏌ц箛姘兼綈鐎规洖顦甸弻鏇熺箾閸喖濮曢梺璇茬箣閻掞妇鎹㈠┑鍡忔灁闁割煈鍠楅悘鎾绘⒑鏉炴壆顦︽い顓犲厴閻涱噣宕�?鑺ユ闂佺粯枪鐏忔瑩藝閵娿儺娓婚柕鍫濇閳锋帡鏌￠崪浣镐喊鐎规洏鍨藉畷锟犳倷閳哄�?�鏉搁梻浣虹帛椤洨鍒掗姘ｆ鐟滃孩绌辨繝鍥舵晝闁挎繂瀛╅悿浣割渻閵堝啫鐏俊顐㈠暣閵嗕線寮崼婵嬪敹闂佺粯鏌ㄩ幖顐︾嵁閸儲鈷掑ù锝囨�?椤曟粎绱掔拠璇ф嫹?閿熶粙鐛繝鍥х疀妞ゆ柨澧介悡瀣攽閻愬弶鈻曞ù婊勭箞閺佹捇鏁撻敓锟??????闂佽鍑界紞鍡涘礈濞戙垺鏅柣鏂垮悑閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曞礈瑜忕壕濂告煕濞嗗浚妲归柕鍥ㄧ箘閳ь剚顔栭崰妤勩亹閸愵喖鐓橀柟杈剧畱闁卞洭鏌曡箛瀣仼缂佺姷鏁诲缁樻媴閸涘﹥鍎撻梺鍝ュ櫏閸嬪﹪骞冭缁绘繈宕堕妸銉ょ暗婵犵數鍋為崹鍫曞春閸愵喖纾婚柟鎹愵嚙�???鍌氼熆鐠虹尨姊楀瑙勬礋濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犻弶鍫㈠亾閿燂拷??闂佽法鍠曟慨銈吤洪幋�???�???闁告劕妯婇崵鏇灻归悩宸剾闁轰礁娲弻锝呂熼崹顔炬闂侀潧鐗炵粻鎾愁潖缂佹ɑ濯村�?�姘煎灡閺侇垶姊虹憴鍕仧濞存粎鍋熼崚鎺撶節濮橆剛顓洪梺缁樏敓�????缂佹顦埞鎴︽倷閺夋垹浠ч梺鎼炲妽濡炰粙宕哄☉銏犵婵°�?�鑳堕崢鍗烆渻閵堝棗濮傞柛濠冩礋瀵悂寮�?崼鐔哄帗濡炪倖鐗楃粙鎺旂矆閸愵喗鐓忛柛銉戝喚浼冮悗娈垮櫘閸撶喎鐣疯ぐ鎺濇晪闁告侗鍓涘Λ顖滅磽閸屾熬�????閿熶粙鎳楅崜浣稿灊妞ゆ牗绮嶅畷鏌ユ煕閺囥劌鐏犵紒鎰殔閳规垿鎮╅煫顓℃姉闂佺粯妫�?鏍惞閸︻厾锛滃┑鈽嗗灥閸嬫劖鏅ラ梻鍌氾拷?锟介崐鎼佸磹閻戣姤鏅搁柨鐕傛�???濠碉紕鍋戦崐鏍垂閻㈢ǹ绠犳慨妞诲亾闁绘侗鍠楃换婵嬪磼閵堝棗缂撻梻渚婃�??閿熻棄鑻晶顔姐亜閺囶亞绉い銏℃礋閺佹捇鏁撻敓�?????缂備讲鍋撻柛鎰ㄦ杺娴滄粓鏌￠崘顭掓嫹?閿熶粙骞忛埄鍐闁绘挸鍑介煬顒佹叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚倷鑳堕�?�濠傗枍閺囥垹绠查柛銉墰�?�撲焦淇婇妶鍛櫣闁告濞婇弻鏇＄疀婵犲喛锟???閿熶粙鏌熼柨瀣仢婵﹥妞藉畷銊︾節閸曨厾鏆ら梺璇插閸戝綊宕ｉ崘銊ф殾闁圭儤顨呮儫闂佸啿鎼崐濠氬储闁秵鈷戦梻鍫熻儐瑜版帒纾匡�??锟芥洖娲ㄩ惌鎾寸箾�?�割喕绨奸柣鎾寸洴閹﹢鎮欓悽鍨啒闂佺ǹ瀛╁Λ鎴﹀箯閿燂拷??闂佽法鍠曟慨銈吤洪弽顓熷亯闁稿繘妫跨换鍡樻叏濠靛棛鐒炬俊鏌ョ畺濮婄儤瀵煎▎鎴犳殸闂佺粯顨嗛幐鎼侊綖韫囨梻�???婵﹩鍓涢敍婊冣攽椤旂煫顏勭暦椤掑嫭鏅搁柨鐕傛嫹?缂傚倸鍊搁崐椋庣矆閿燂拷?椤㈡牠宕卞▎鎰闂佺粯鍔欏褔宕瑰┑鍡忔斀闁绘ê寮堕幖鎰版煟閹惧娲撮柡灞剧〒娴狅箓宕滆閸ｎ喚绱撴担鍝勑ｉ柤褰掔畺閳ユ棃宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣绮欓崠鈩冩暰濠电偛寮堕…鍥╁垝鐎ｎ喖绠抽柟瀛樻煥閻楁岸姊洪崨濠冪５闁哄懏鐟ч懞杈╂嫚瀹割喗�?�岄梺闈涚墕閹虫劗绮绘导瀛橈�??锟芥慨妯煎帶婢ц揪�????閿熺瓔鍠楁繛濠囧极閹版澘宸濇い蹇撴噺閺夋悂姊绘担鍝勪缓闁稿氦浜竟鏇㈩敇閵忕姵锟??????闂備礁鎼ú锕傛晪婵犳鍠栭崐褰掑Φ閸曨垰顫呴柨娑樺閿燂拷??闂備胶顢婇崑鎰偘閵夆晛�?堟繝闈涱儏濮瑰弶銇勮箛鎾跺闁抽攱甯￠弫鎾绘晸閿燂拷??????闂傚倷鑳堕崢褔宕幐搴㈡珷閹兼番鍔岀粈鍡涙煙閻戞﹩娈㈤柡浣哥Ч閺岋綁骞囬鐔虹▏婵炲瓨绮撴禍璺侯潖濞差亜浼犻柛鏇ㄥ墮閸嬪秹姊洪幖鐐插闁硅櫕鎸哥叅闁秆勵殕閳锋帒霉閿濆懏鎲哥紒澶屽劋娣囧﹪顢曢�?鈥充淮闂佽鍠氶崑銈夊极閸愵喖纾兼慨妯诲敾缁辫鲸绻濆▓鍨灍闁靛洦鐩畷鎴﹀箻缂佹鍘搁柣蹇曞仩椤曆勬叏閸岀偞鐓欐い鏂挎惈閳ь剚绻傞悾鐑藉箳閹存梹�???????闂傚倸鍊峰ù鍥敋瑜忛�?顒佺▓閺呯娀銆佸▎鎾冲唨妞ゆ挾鍋熼悰銉╂⒑閸濆嫭宸濆┑顔芥尦瀹曠懓鈹戦崶鈺冾啎闂佺硶鍓濋敋濠殿喖鍟扮槐鎺�?嫚閸欏妫﹂梺鍝勭灱閸犳牕顫忛懡銈傚亾閻㈢櫥瑙勪繆娴犲鈷戦柛婵嗗閸ｈ櫣绱掗鑺ュ磳鐎殿喛顕ч埥澶愬閻樻鍟岄梻浣告啞閸旓附绂嶅▎鎾存優閹兼番鍔嶉埛鎴︽⒒閸喓銆掑褎娲�?妵鍕晜閸喖绁�?梺绯曟櫆閻╊垶鐛�?幒锟??绠犻柕濞垮劤缁夋椽鏌℃担鐟板鐎规洖銈搁幃銈嗘媴瀹勭増鎲㈤梻鍌欑劍閻綊宕洪崟顖氬�?�闂侇剙绉甸崕搴€亜閺嶎偄浠滈柦鍐枑缁绘盯骞嬪▎蹇曚患缂備緡鍋勭粔褰掑蓟閻旂厧绠氱憸宥夛拷?锟介幎鑺ョ厸闁糕剝鍔曢埀顒佺箞楠炲啫螖閸愨晛鏋傞梺鍛婃处閸撴盯藝閵娧呯＝濞撴艾娲ら弸娑㈡煟椤撶儑�????閿熻棄鐣峰ú顏勵潊闁斥晛鍟崝鍛存⒑闂堟胆褰掑磿閹剁瓔鏁婇柟鍓х帛閳锋垿鏌涘☉姗堝伐濠殿喒鍋撻梻浣告惈閹冲繒鍒掑畝鍕厺鐎广儱顦獮銏＄箾閹寸偟鎲块柟椋庣帛缁绘稒娼忛崜褏袣婵犳鍠撻崐�???鈽夐悽绋块唶闁哄洨鍠撻崢閬嶆⒑閹稿海绠撶紒缁樺浮閹箖宕归顐ｎ啍闂佺粯鍔樼亸娆戠不婵犳碍鐓涘ù锝堫潐瀹曞矂鏌ㄩ悤鍌涘�????
        .bid(bid),      
        .bresp(bresp),    
        .bvalid(bvalid),        
        .bready(bready)         
    );

    cache_AXI u_cache_AXI(
        .clk(aclk),
        .rst(rst),    // low active

    //icache read
        .inst_ren_i(icache_ren),
        .inst_araddr_i(icache_araddr),
        .inst_rvalid_o(icache_rvalid),
        .inst_rdata_o(icache_rdata),
        .icache_ren_received(icache_ren_received),
        .icache_flush_flag_valid(icache_flush_flag_valid),

    //dcache read
        .data_ren_i(dcache_ren),
        .data_araddr_i(dcache_araddr),
        .data_rvalid_o(dcache_rvalid),
        .data_rdata_o(dcache_axi_data_block),
        .dcache_ren_received(dcache_ren_received),

    //dcache write
        .data_wen_i(dcache_wen),
        .data_wdata_i(dcache_wdata),
        .data_awaddr_i(dcache_awaddr),
        .data_bvalid_o(dcache_bvalid),

        .cache_axi_write_pre_ready(cache_axi_write_pre_ready),

    //ready to cache
        .dev_rrdy_o(dev_rrdy_to_cache),
        .dev_wrdy_o(dev_wrdy_to_cache),
    //uncache to icache
        .iuncache_ren_i(iuncache_ren),
        .iuncache_raddr_i(iuncache_raddr),
        .iuncache_rvalid_o(iuncache_rvalid),
        .iuncache_rdata_o(iuncache_rdata), 

    //uncache to dcache
        .duncache_ren_i(duncache_ren),
        .duncache_raddr_i(duncache_raddr),
        .duncache_rvalid_o(duncache_rvalid),
        .duncache_rdata_o(duncache_rdata),

        .duncache_wen_i(duncache_wen),
        .duncache_wstrb(duncache_wstrb),
        .duncache_wdata_i(duncache_wdata),
        .duncache_waddr_i(duncache_waddr),
        .duncache_write_resp(duncache_write_finish),

    //AXI communicate
        .axi_ce_o(axi_ce_o),
        .axi_wsel_o(axi_wsel),   // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁绘劦鍓欓崝銈囩磽�?�ュ拑韬拷?锟筋喖顭烽幃銏ゅ礂鐏忔牗瀚介梺璇查叄濞佳勭珶婵犲伣锝夘敊閸撗咃紲闂佺粯鍔﹂崜娆撳礉閵堝鏅搁柨鐕傛嫹?闂備緡鍓欑粔鎾倿閸偁浜滈柟鐑樺灥閳ь剙缍婇弫鎾绘晸閿燂�???闂備浇顕э�??锟解晠宕欒ぐ鎺戠煑闁告劑鍔庨弳锔兼嫹?閿熻姤娲栧ú銈壦夊鑸碉拷?锟介柨婵嗗暙婵＄儤鎱ㄧ憴鍕垫疁婵﹥妞藉畷鐑筋敇閻愭彃顬嗛梻浣规偠閸斿瞼绱炴繝鍌滄殾闁规壆澧楅崐鐑芥煟閹寸伝顏呯椤撶偐�?介柣妯款嚋�?�搞儵鏌ㄩ悤鍌涘�????闂備浇顕э�??锟解晠顢欓弽顓炵獥婵°倕鎳庣粻鏍煕鐏炴儳鍤柛銈嗘礀闇夐柣妯烘▕閸庢盯鏌℃担鍛婂枠闁哄矉缍佸顒勫箰鎼淬垹鍓垫俊銈囧Х閸嬬偤宕濆▎蹇ｆ綎缂備焦蓱婵挳鎮峰▎蹇擃仼濞寸姭鏅犲铏圭矙閸喚妲伴梺鎼炲姀濞夋盯鎮鹃悜钘夊嵆闁靛骏绱曢崝鍫曟煥閻曞倹锟???????闂傚倸鍊风粈�???宕崸锟??绠规い鎰剁畱閻ゎ噣鏌熷▓鍨灈妞ゃ儲鑹鹃埞鎴�?磼濮橆厼鏆堥梺缁樻尰閻熲晛顫忛敓�???????闁诲孩顔栭崰姘跺磻閹捐埖宕叉繛鎴欏灩闁卞洭鏌ｉ弮鍥仩闁绘挸顦甸弫鎾绘晸閿燂�???????闂備椒绱徊鍓ф崲閸儲鏅搁柨鐕傛�??婵＄偑鍊栫敮鎺炴�??閿熺瓔鍓涚划锝呂旈崨顔惧幐閻庡箍鍎辨鎼佺嵁閺嶎偆纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍓涢幑鍕Ω閿旂瓔鍟庢繝鐢靛█濞佳囧磹閹间礁绠熼柨鐔哄Т绾惧鏌涢弴銊ョ仭闁绘挻娲樼换婵嬫濞戞瑯妫炲銈呯箚閺呮粎鎹㈠☉銏犻唶婵炴垶锚婵箑鈹戦纭峰伐妞ゎ厼鍢查悾鐑藉箳閹存梹鐎婚梺瑙勬儗閸橈�??锟解叺闂傚�?�鍊烽懗鍫曪�??锟芥繝鍥舵晪婵犲﹤鎳忓畷鍙夌�?闂堟稒顥犻柡鍡畵閺屾盯鏁傜拠鎻掔闂佸摜濮村Λ婵嬪蓟閿燂�?????闁诲孩顔栭崰鏍ь焽閳ユ剚娼栨繛宸簻閹硅埖銇勯幘顖氬⒉妞ゅ孩顨婂娲传閵夈儛锝夋煟濡ゅ啫鈻堟鐐插暣閸ㄩ箖骞囨担鐟扮紦闂備緤�????閿熻棄鑻晶杈炬�??閿熺瓔鍠栭�?�鐑藉箖閵忋倕宸濆┑鐘插鑲栨繝寰峰府锟???閿熺晫寰婃禒瀣柈妞ゆ牜鍎愰弫渚婃嫹?閿熷鍎遍ˇ浼村煕閹寸姷纾奸悗锝庡亽閸庛儵鏌涙惔銏犲闁哄本鐩弫鎾绘晸閿燂拷??闂佽崵鍟块弲鐘绘偘閿燂拷?瀹曟﹢濡告惔銏☆棃鐎规洏鍔戦、锟??鎮㈡搴涘仩婵犵绱曢崑鎴﹀磹閺嶎厼绠板Δ锝呭暙绾捐銇勯幇鍓佺暠妞ゎ偄鎳�?獮鎺楁惞椤愩値娲稿┑鐘诧工閻�?﹪鎮¤箛鎿冪唵闁煎摜鏁搁埥澶嬨亜閳哄﹤澧扮紒杈ㄥ浮閹晠骞囨担鍝勫Ш缂傚倷娴囨ご鍝ユ暜閿燂拷?椤洩绠涘☉妯溾晠鏌ㄩ悤鍌涘�??闂傚倸顦粔鐟邦潖濞差亝鍋￠柡澶嬪浜涢梻浣侯攰濞呮洟鏁嬮梺浼欑悼閸忔﹢銆侀弴銏℃櫢闁跨噦锟???缂備讲鍋撻悗锝庡墰濡垶鏌ｉ敓锟???閻擃偊顢旈崨顖ｆ�?????闂備緤锟???閿熻棄鑻晶杈炬�??閿熻姤娲滈崰鏍�??锟藉Δ鍛＜婵﹩鍓涢悿鍕⒒閸屾熬锟???閿熺晫娆㈠鑸垫櫢闁跨噦�?????闂傚倷鑳舵灙閻庢稈鏅滅换娑欑�?閸屾粍娈惧┑鐐叉▕娴滄繈寮查弻銉︾厱闁靛鍨抽崚鏉棵瑰⿰鍛壕缂佺粯鐩畷鐓庘攽閸粏妾搁梻浣告惈椤戝棛绮欓幒锟??桅闁告洦鍨奸弫鍥煟濡绲绘鐐差儔閹鈻撻崹顔界彯闂佺ǹ顑呴敃顏堟偘閿燂�??瀹曞爼顢楁径瀣珝闂備胶绮崝妤呭极閹间焦鍋樻い鏂跨毞锟??浠嬫煟濡櫣浠涢柡鍡忔櫅閳规垿顢欑喊鍗炴�??濠殿喗锚瀹曨剟宕拷?锟界硶鍋撶憴鍕８闁稿酣娼ч悾鐑斤�??锟介幒鎾愁伓?闂佽法鍠曟慨銈堝綔闂佸綊顥撶划顖滄崲濞戞瑦缍囬柛鎾楀嫬浠归梻浣侯攰濞呮洟骞戦崶顒婃嫹?閿熻棄顫濋钘夌墯闂佸憡渚楅崹鎶芥晬濠婂牊鐓熼柣妯哄级婢跺嫮鎲搁弶鍨殻闁糕斁鍋撻梺璺ㄥ櫐閿燂拷??濠电偟銆嬬换婵嬪箖娴兼惌鏁婇柦妯侯槺缁愮偞绻濋悽闈涗户闁稿鎹囬敐鐐差吋婢跺鎷洪梻鍌氱墛缁嬫挾绮婚崘娴嬫斀妞ゆ梹鍎抽崢瀛樸亜閵忥紕鎳囨鐐村浮瀵噣宕掑⿰鎰棷闂傚�?�鑳舵灙闁哄牜鍓熼幃鐤樄鐎规洘绻傞濂稿幢閹邦亞鐩庢俊鐐�??锟介幐楣冨磻閻愬搫绐楁慨�???鐗婇敓锟????闂佽法鍠曟慨銈吤鸿箛娑樺瀭濞寸姴顑囧畵锟??鏌�?�鍐ㄥ濠殿垱鎸抽弻娑滅疀閹垮啯效闁诲孩鑹鹃妶绋款潖缂佹ɑ濯撮柛娑橈工閺嗗牏绱撴担鍓插剱闁搞劌娼″顐﹀礃椤旇姤娅滈梺鎼炲労閻撳牓宕戦妸鈺傗拻濞撴艾娲ゆ晶顔剧磼婢跺本鏆柟顕嗙�?瀵挳锟??閿涘嫬骞楁繝纰樻閸ㄧ敻顢氳閺呭爼顢涘☉姘鳖啎闂佸壊鍋嗛崰鎾绘儗锟??鍕厓鐟滄粓宕滃┑�?�剁稏濠㈣泛鈯曞ú顏呮櫢闁跨噦�????閻庤娲樼换鍌炲煝鎼淬劌绠婚悹楦挎閵堬箓姊绘担瑙勫仩闁稿孩妞藉畷婊冾潩鐠鸿櫣锛涢柣搴秵閸犳鎮￠弴鐔翠簻闁归偊鍠栧瓭闂佽绻嗛弲婊堬�??锟介妷鈺傦拷?锟介柡澶嬪灥椤帒鈹戦纭烽練婵炲拑缍侀獮鎴�?礋椤栨鈺呮煏婢舵稑顩憸鐗堝哺濮婄粯鎷呴悜妯烘畬闂佽法鍣﹂敓锟???????闂傚倸鍊搁崐宄懊归崶顒夋晪鐟滄柨鐣峰▎鎾村仼閿燂�??閳ь剛绮堟繝鍥ㄧ厱闁斥晛鍟伴埥澶岀磼閳ь剟宕奸悢铏诡啎闂佺懓鐡ㄩ悷銉╂�?�椤忓牊鐓曢幖绮规闊剟鏌＄仦鍓ф创妞ゃ垺娲熼幃鈺呭箵閹烘埈娼ラ梻鍌欒兌鏋柨鏇畵瀵偅绻濆顒傜暫閻庣懓瀚竟�?�几鎼淬劎鍙撻柛銉ｅ妽閹嫬霉閻樻彃鈷旂紒杈ㄦ尰閹峰懘骞撻幒宥咁棜闂傚倷绀�?幉锟犲礉閿曞倸绐楁俊銈呮噹绾惧鏌曟繝蹇氱濞存粍绮撻弻鈥愁吋閸愩劌顬嬮梺�?�犳椤︽壆鎹㈠☉銏犵妞ゆ挾鍋為悵婵嬫⒑閸濆嫯顫﹂柛鏂跨焸閸╃偤骞嬮敓�????闁卞洦绻濋棃娑欏櫧闁硅娲樻穱濠囧Χ閸�?晜顓规繛瀛樼矋閻熲晛鐣烽敓鐘茬闁肩⒈鍓氬▓楣冩⒑缂佹ɑ灏紒銊ョ埣�?�劍绂掞拷?锟筋偓锟???閿熶粙鏌ㄥ┑鍡欏嚬缂併劌銈搁弻锟犲幢閿燂�??闁垱鎱ㄦ繝鍌ょ吋鐎规洘甯掗埢搴ㄥ箳閹存繂鑵愮紓鍌氾�??锟界欢锟犲闯閿燂�??瀹曞湱鎹勬笟顖氭婵犵數濮甸懝鐐�?劔闂備礁纾幊鎾惰姳闁秴纾婚柟鎹愵嚙锟??鍐煃閸濆嫸�????閿熶粙宕濋崨瀛樷拺闂傚牊绋堟惔鐑芥⒒閸曨偄顏╅柍璇茬Ч閿燂�??闁靛牆妫岄幏娲煟閻樺厖鑸柛鏂胯嫰閳诲秹骞囬悧鍫㈠�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉绻濋弫鎾绘晸閿燂�???闂佸摜濮甸悧鐘荤嵁閸愵収妯勯悗瑙勬礀閵堟悂骞冮姀銈呬紶闁告洦鍋呴濂告⒒閸屾熬锟???閿熺晫绮堥敓�????楠炲鏁撻悩鎻掞�??锟介柣鐔哥懃鐎氼參宕ｈ箛娑欑厵缂備降鍨归弸娑㈡煟閹捐揪鑰块柡�???鍠愬蹇斻偅閸愨晪锟???閿熶粙姊虹粙娆惧剱闁告梹鐟╅獮鍐ㄎ旈崨顓熷祶濡炪倖鎸鹃崐顐﹀鎺虫禍婊堟煏婢舵稑顩紒鐘愁焽缁辨帗娼忛妸�???闉嶉梺鐟板槻閹虫ê鐣烽敓锟???????闂傚倸鍊烽悞锕傚箖閸洖�?夐敓�????閸曨剙浜梺缁樻尭鐎垫帡宕甸弴鐐╂斀闁绘ê鐤囨竟锟??骞嗛悢鍏尖拺闁告劕寮堕幆鍫ユ煕婵犲�?�鍟炵紒鍌氱Ч閹瑩鎮滃Ο閿嬪缂傚倷绀�?鍡嫹?閿熺獤鍐匡拷?锟介柟娈垮枤绾惧ジ鎮楅敐搴�?�簻闁诲繐鐡ㄩ妵鍕閳╁喚妫冮梺璺ㄥ櫐閿燂�?????闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鎯у⒔濞呫垽骞忛敓�?????闂佽法鍠曞Λ鍕舵嫹?閿熺瓔鍙冨畷宕囧鐎ｃ劋姹楅梺鍦劋閸ㄥ綊宕愰悙鐑樺仭婵犲﹤鍠氶敓锟???閻庢鍠楅幃鍌氼嚕娴犲鏁囬柣鏂挎惈楠炴劙姊绘担瑙勫仩闁稿寒鍨跺畷鏇㈡焼瀹ュ棴锟???閿熶粙鏌嶉崫鍕殶缁炬儳銈搁弻鐔兼焽閿燂�??瀵偓绻涢崼鐔虹煉闁哄矉�????閿熺晫鏆嗛悗锝庡墰閻�?牓鎮楃憴鍕闁绘牕銈稿畷娲焺閸愨晛顎撻梺鍦帛鐢﹥绔熼弴銏�?拺闁圭ǹ娴风粻鎾绘煙閸愬樊妲搁崡閬嶆煕椤愮姴鍔滈柣鎾崇箻閻擃偊宕堕妸锔绢槬闁哥喓枪椤啴濡惰箛娑欙�??锟藉┑鐘灪閿曘垽鍨鹃弮鍫濈妞ゆ柨妲堣閺屾盯鍩勯崗锟??浜鍐参旀担铏圭槇濠电偛鐗嗛悘婵嬪几閵堝鐓曢煫鍥ㄦ�?�閻熸嫈娑㈡偄婵傚瀵岄梺闈涚墕濡稒鏅堕鍌滅＜閻庯綆鍋呯亸纰夋嫹?閿熺瓔鍟崶褏鍔�?銈嗗笒鐎氼參鍩涢幋鐐村弿闁荤喓澧楅幖鎰版煟韫囨挸绾х紒缁樼⊕閹峰懘宕�?幓鎺撴闂佺懓顫曢崕閬嶅煘閹达附鍋愰柛顭戝亝濮ｅ嫰姊虹粙娆惧剱闁烩晩鍨堕獮鍡涘炊閵娿儺鍤ら梺鍝勵槹閸ㄥ綊鏁嶅▎蹇婃斀闁绘绮☉褎銇勯幋婵囧櫧缂侇喖顭烽、娑㈡�?�鐎电ǹ骞嶉梺鍝勵槸閻楁挾绮婚弽褜鐎舵い鏇�?亾闁哄本绋撻�?顒婄秵娴滄粓顢旈銏＄厸閻忕偛澧介�?�鑲╃磼閻樺磭鈽夋い顐ｇ箞椤㈡牠骞愭惔锝嗙稁闂傚倸鍊风粈�???骞夐敓鐘虫櫇闁冲搫鍊婚�?�鍙夌節闂堟稓澧涳拷?锟芥洖寮剁换婵嬫濞戝崬鍓遍梺绋款儍閸旀垵顫忔繝姘唶闁绘棁�???濡晠姊洪悷閭﹀殶闁稿繑锚椤繘鎼归崷顓犵厯濠电偛妫欓崕鎶藉礈闁�?秵鈷戦柣鐔哄閸熺偤鏌熼纭锋嫹?閿熻棄鐣峰ú顏勵潊闁绘瑢鍋撻柛姘儏椤法鎹勯悮鏉戜紣闂佸吋婢�?悘婵嬪煘閹达附鍊烽柡澶嬪灩娴犳悂姊洪懡銈呮殌闁搞儜鍐ㄤ憾闂傚倷绶￠崜娆戠矓閻㈠憡鍋傞柣鏃傚帶缁犲綊鏌熺喊鍗炲箹闁诲骏绲跨槐鎺撳緞閹邦厽閿梻鍥ь槹缁绘繃绻濋崒姘间紑闂佹椿鍘界敮妤呭Φ閸曨垰顫呴柍鈺佸枤濡啫顪冮妶鍐ㄧ仾闁挎洏鍨介弫鎾绘晸閿燂�???闂備焦�?�х粙鎴�??閿熺瓔鍓熼悰�???骞囬悧鍫氭嫼闁荤姴娲╃亸娆戠不閹惰姤鐓曢悗锝庡亞閳洟鏌￠崨鏉跨厫缂佸�?�甯為埀顒婄秵娴滅偤宕ｉ�?�???鈹戦悩顔肩伇闁糕晜鐗犲畷婵嬪�?椤撶喎浜楅梺鍛婂姦閸犳鎮￠�?鈥茬箚妞ゆ牗鐟ㄩ鐔镐繆椤栨氨澧涘ǎ鍥э躬楠炴捇骞掗幘铏畼闂備線娼уú銈忔�??閿熸垝鍗抽妴�???寮撮�?鈩冩珳闂佹悶鍎弲婵嬪储濠婂牊鐓熼幖娣�??锟藉鎰箾閸欏鐭掞拷?锟芥洏鍨奸ˇ褰掓煕閳哄啫浠辨鐐差儔閺佹捇鏁撻敓锟????濡ょ姷鍋戦崹浠嬪蓟�?�ュ浼犻柛鏇�?�煐閿燂�???闂佽法鍠撻弲顐ゅ垝婵犲浂鏁婇柣锝呯灱閻﹀牓姊哄Ч鍥х伈婵炰匠鍐╂瘎闂傚�?�娴囧銊╂倿閿曞�?�绠栭柛灞炬皑閺嗭箓鏌燂�??锟芥濡囨俊鎻掔墦閺屾洝绠涙繝鍐╃彆闂佸搫鎷嬫禍婊堬�??锟介崘顔嘉ч柛鈩兠拕濂告⒑閹肩偛濡肩紓宥咃工閻ｇ兘骞掗敓�????鎯熼悷婊冮叄瀹曚即骞囬鐘电槇闂傚�?�鐗婃笟妤呭磿韫囨洜纾奸柣娆屽亾闁搞劌鐖煎濠氬Ω閳哄倸浜為梺绋挎湰缁嬫垿顢旈敓锟????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ら娑㈡⒑缂佹ɑ鐓ユ俊顐ｇ懇楠炲牓濡搁妷顔藉瘜闁荤姴娲╁鎾寸珶閺囥垺鈷掑ù锝囨嚀椤曟粎绱掔拠鎻掝伃鐎规洘鍨块幃鈺呮偨閸忓摜鐟濇繝鐢靛仦閸垶宕归悷鎷�?稑顫滈埀顒勫箖瑜版帒鐐婃い蹇撳婢跺嫰姊洪崫銉バ㈤柨鏇ㄤ簻椤繐煤椤忓懎娈ラ梺闈涚墕閹冲繘鎮�?ú顏呪拻闁稿本鑹鹃鈺冪磼婢跺本锟??闁伙絿鍏�?獮鍥�?级鐠侯煈鍟嬮梻浣哥秺濞佳囨�?�閺囥垹�?傞柣鎰靛墯椤ュ牞�????閿熻姤娲忛崝鎴︼�??锟藉▎鎴炲枂闁告洦鍋掓导鏍⒒閸屾熬�????閿熺晫娆㈠顒夌劷濞村吋鐟﹂敓锟????闂佽法鍠曞Λ鍕儗閸屾氨鏆﹂柕蹇ョ磿闂勫嫮绱掞�??锟筋厽纭舵い锔诲櫍閺岋絾鎯旈婊呅ｉ梺鍛婃尰缁嬫挻绔熼弴鐔洪檮闁告稑锕ゆ禒顖炴⒑閹肩偛鍔�?柛鏂跨灱瀵板﹥绻濆顓犲幐闂佺硶妲呴崢鍓х矓閿燂拷?閺岀喓绮欓崠陇鍚梺璇�?�枔閸ㄨ棄鐣峰Δ鍛殐闁宠桨绀佺粻浼存⒑鐠囨煡顎楃紒鐘茬Ч�?�曟洘娼忛�?�鎴烆啍闂佸綊妫块懗璺虹暤娴ｏ拷?锟界箚闁靛牆鎳忛崳娲煟閹惧啿鏆ｆ慨濠冩そ�?�曞綊顢氶崨顓炲闂備浇顕х换鍡涘疾濠靛牊顫曢柟鐑樻尰缂嶅洭鏌曟繛鍨姢妞ゆ垵鍊垮娲焻閻愯尪�?�板褍澧界槐鎾愁吋閸涱噮妫﹂悗瑙勬磸閸ㄤ粙骞冮崜褌娌柟顖嗗啫绠查梻鍌欑閹诧繝骞愰悜鑺ュ殑闁告挷�?�?ˉ姘攽閸屾碍鍟為柣鎾跺枑娣囧﹪顢涘┑鍥朵哗闂佹寧绋戠粔褰掑蓟濞戞ǚ鏋庨悘鐐村灊婢规洟姊婚崒姘炬�??閿熺晫绮堥敓�????楠炴牠顢曢妶鍡椾粡濡炪�?�鍔х粻鎴犵矆婢舵劖鐓欓悗娑欘焽缁犮儵鏌涢妶鍡樼闁哄备鍓濆鍕舵�??閿熺瓔浜濋鏇㈡⒑缂佹ɑ鐓ラ柛姘儔楠炲棝鎮欓悜妯锋嫼濡炪倖鍔х徊鍧�?�?閺囥垺鐓曢悗锝庝簼閸ｅ綊鏌嶇憴鍕伌闁轰礁绉瑰畷鐔碱敃閳╁啯绶氶梻鍌欒兌鏋柨鏇樺劦閹囧即閻樻彃鐤鹃梻鍌欑閸熷潡骞栭锟??鐤柟娈垮枤閻棗鈹戦悩鎻掍喊闁瑰嚖�????闂佽法鍠曞Λ鍕綖濠靛鏅查柛娑卞墮椤ユ岸姊婚崒娆戠獢婵炰匠鍏炬盯寮崒娑卞仺濠殿喗锕╅崜锕傚吹閺囥垺鐓欑紓浣靛灩閺嬫稒銇勯銏�?�殗闁哄苯绉归崺鈩冩媴閸涘﹥顔夐梻浣虹帛缁诲啴鎮ч悩缁樻櫢闁跨噦锟?????闂備緤锟???閿熻棄鑻晶浼存煕鐎ｎ偆娲撮柟宕囧枛椤㈡稑鈽夊▎鎰娇闂備浇顫夐鏍窗濮樺崬顥氶柛蹇曨儠娴滄粓鏌￠崒姘变虎闁抽攱妫冮幃浠嬵敍濞戞熬�????閿熺晫绱掓潏銊ョ缂佽鲸甯掕灒闁兼祴鏅濋弳銈嗕繆閻愵亷锟???閿熶粙宕戦崨顖涘床闁割偁鍎�?顑跨窔閺佹捇鏁撻敓锟????闂佽鍠掗弲鐘荤嵁閹捐绠抽柡鍐拷?锟藉鏍⒒閸屾熬锟???閿熶粙宕愰幖浣哥９鐎瑰嫭鍣磋ぐ鎺戠�?�妞ゆ帒锕︾粙蹇旂節閵忥絾纭鹃柨鏇畵�?�娊鏁傞幋鎺旂畾濡炪�?�鐗滈崑鐐烘晬閻斿吋鐓熼柟鐑樺煀�???鑽ょ磼缂佹娲达�??锟芥洖宕灒閻犲洤妯婃导鍥⒒娴ｈ鍋犻柛搴㈡そ瀹曟粌顫濈捄铏规煣濠电姴锕ら悧濠囨偂閺囥垻鍙撻柛銉ｅ妽閿燂拷?闁汇埄鍨甸崺鏍Φ閿燂�?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殜閺岋繝宕堕埡浣癸拷?锟介梺鍛婄懃缁绘﹢寮婚弴銏犻唶婵犻潧娲ゆ禒鐐繆閵堝繒鐣虫繛澶嬫礋閺佹捇鏁撻敓锟????濠电姷鏁搁崑鐐哄垂閸洩�????閿熶粙宕堕浣规珫闂佺粯鏌ㄩ崥�?�煕閹烘埊�????閿熻棄顫濋浣规倷婵犫拃灞芥灓缂佽鲸甯楀鍕熼悜妯煎綆??濠碉紕鍋戦崐鏍暜婵犲洦鍊块柨鏇炰紪閿燂�??????闂備礁鎼ú銊╁闯閿曞倹锟??闁圭ǹ绨烘禍婊堟煏韫囥儳纾块柟鍐叉川閳ь剝顫夊ú鏍ь嚕閸撲胶鍗氶柣鏃傗拡閺佸秵鎱ㄥ鍡楀箹妞わ腹鏅犲铏圭磼濡闉嶅┑鐐跺皺閸犳牕顕ｇ拠宸悑濠㈣泛锕﹂崢鍛婄箾鏉堝墽鎮奸弸顏嗙磼閻樹警鍤欐い顏勫暣婵″爼宕ㄩ婊庡敹闂備胶绮�?�鍛涘Δ浣规珡闂備礁鎲￠悷銉┧囬鐐�?床闁糕剝绋掗悡蹇涙煕椤愶絿绠撴い蹇ｅ墴閺屾稖绠涢幘鍓佷紘缂備浇椴哥敮锟犲春閿燂拷??闂備胶枪椤戝棝骞愰懡銈嗗床婵犻潧顑嗛崑銊╂⒒閸喓鈼ョ紒顔肩埣濮婅櫣绱掑鍡樼暥濠碘槅鍋呯换鍫ョ嵁閸愩剮鐔烘偘閳╁啯鏉搁梺璺ㄥ櫐閿燂�???????闂佽法鍣﹂敓�????????缂傚倷绀�?ˇ閬嶅极婵犳艾绠栭柨鐔哄Т閸楁娊鏌ｉ弮鍥仩妞ゆ梹娲熷铏瑰寲閺囩偛鈷夊銈冨妼閻楀繒鍒掔紒妯侯嚤閻庢稒顭囬崢鎼佹⒑缁洖澧叉い顓炴喘楠炲﹪宕熼娑氬帾闂佹悶鍎滈崘鍙ョ磾闁诲孩顔栭崰妤呭箰閹舵枻锟???閿熶粙寮�?崼婵嗭拷?锟藉┑鐐叉噽閸庛倗鍒掗幘璇茬畺婵°倕鍟崰鍡涙煕閺囥劌澧版い锔哄姂濮婃椽骞愭惔鈥虫懙濠碘槅鍋傞悞锟??顕ラ崟顖氱疀妞ゆ挶鍔嶉敓�?????闂佽法鍠嶇划娆撳蓟閵娿儮�?介柛鈩冪懃閸ゎ剛绱撴担闈涘婵☆偄�?�伴垾锕傛嚄椤栵絾顎囬梻浣规偠閸斿繐鈻斿☉顫稏闊洦娲滅壕鍏间繆椤栨繍鍤欐い搴㈡尵缁辨挻鎷呴崜鎻掑壉濡炪�?�鍨堕悷銉ㄧ亱閻庡厜鍋撻柛鏇ㄥ厴閹疯櫣绱撴担鍓插剱妞ゆ垶鐟╁畷鏇＄疀閺傚墽绠氬銈嗗姧缁茶法绮婚幘缁樼厽闁挎繂顦伴弫閬嶆倵闂堟稏鍋�??锟筋喖鐖奸獮瀣偑閳ь剟宕拷?锟筋喗鈷戦柤濮愶�??锟藉瓭濠电偠顕滅粻鎺�?Φ閹版澘绀冩い鏃囧亹閿涙盯鎮楅獮鍨姎妞わ缚鍗抽崺娑㈠箣閿旂晫鍘遍梺鐟板⒔閹虫捇鎯冨ú顏呯厱婵☆垵宕靛ú鎾煛鐏炴儳鍠曢柟鍑ゆ�???????闂傚倷鑳堕幊鎾剁不�?�ュ鍨傞柦妯侯槺閺嗭箓鏌涘Δ鍐ㄤ汗婵℃彃鐗婄换娑㈠幢濡櫣浠村Δ鐘靛仦椤ㄥ﹤顫忕紒妯诲闁告縿鍎虫闂備胶枪椤戝懘鏁冮鍕殾婵犲﹤鍠氬鈺呮偣妤︽寧顏犻柛妯绘そ濮婃椽宕崟�???鍋嶉梺鎼炲妽濡炰粙骞冮敓鐘插嵆闁靛繒濮烽鎰版煛婢跺﹦澧曞褏鏅竟鏇犳崉閵娧咃紲闂佺粯锚濡﹪鎮℃總鍛婄厸閿燂�??閳ь剟宕伴弽顓ㄦ嫹?閿熻棄鈻庨幋鐘烩攺闁诲函缍嗛崑鍡涘级閿燂�?????闂備礁鎼ú銊╁磻閻旇櫣鐭撻柣鎴炃滄禍婊堟煏韫囧﹤澧查敓锟???鐎ｎ喗鏅搁柨鐕傛�???闂傚倸鍊革拷?锟筋剙煤椤撱垺鏅搁柨鐕傛�????婵犳鍠栭敃锔惧垝椤栫偛绠柛娑卞灣妞规娊鎮楅敐搴濈凹闁伙絼鍗冲缁樻媴閸涘﹥鍠愭繝娈垮枤閺佸鐛幋锟??鐐婄憸蹇涘汲閿旂偓鍠愰柣�???鐗嗙粭姘舵�?�閻㈤潧孝妞ゎ叀娉曢幑鍕�?�濡粯瀚虫繝鐢靛仜閻楁挾绮婚弽褜娼栨繛宸簻缁犱即骞栨潏鍓у矝婵℃彃鐗撻弻锝嗘償閵忕姴姣堥梺鍝ュУ绾板秶绮嬪澶婄濞达絿鎳撴禒娲⒑濮瑰洤鐏�?柡浣规�?�閺佸秴饪伴崼鐔叉嫼闂傚倸鐗婇懗鍡氥亹閹烘垹锛熷銈嗙墱閸嬫盯鎮為崹顐犱簻闁圭儤鍩婇弨濠氭煥閻曞倹锟???

    //AXI read
        .rdata_i(axi_rdata),
        .rdata_valid_i(axi_rdata_valid),
        .axi_ren_o(axi_ren),
        .axi_rready_o(axi_rready),
        .axi_raddr_o(axi_raddr),
        .axi_rlen_o(axi_rlen),

    //AXI write
        .wdata_resp_i(axi_wdata_resp),  // 闂傚倸鍊搁崐鎼佸磹閹间礁纾归柟闂寸绾惧綊鏌熼梻瀵割槮缁炬儳缍婇弻鐔兼⒒鐎靛壊妲紒鐐劤缂嶅﹪寮婚悢鍏尖拻閻庨潧澹婂Σ顔剧磼閻愵剙鍔ょ紓宥咃躬�?�鎮㈤崗灏栨嫽闁诲酣娼ф竟濠偽ｉ鍓х＜闁诡垎鍐ｆ寖闂佺娅曢幑鍥灳閿燂拷?????婵＄偑鍊曠换鎰板箠韫囨挾鏆﹂柟鎯板Г閳锋垶绻涢懠棰濆殭妤犵偞鐗楁穱濠囶敃閿濆洨鐤勯悗娈垮枛椤攱淇婇幖浣哥厸闁稿本鐭花浠嬫⒒娴ｅ懙褰掑嫉椤掑倻鐭欓柟杈惧瘜閿燂拷???婵犵數濮撮惀澶屾暜椤旇棄�????闂佽法鍠曟慨銈夊箞閵娾晜鍊婚柦妯侯槺閿涙稑鈹戦悙鏉戠亶闁瑰磭鍋ゅ畷鍫曨敆娴ｉ晲缂撶紓鍌欑椤戝棴�????閿熺獤鍥拷?锟芥い鎺戝閳锋垿鏌ｉ悢鍛婄凡闁抽攱姊荤槐鎺楊敋閸涱厾浠搁悗瑙勬礃閸ㄥ潡鐛崶顒佸亱闁割偁鍨归獮妯肩磽娴ｅ搫浜炬繝銏∶悾鐑筋敆娴ｈ鐝风紓鍌欑劍鐪夌紒璇叉閺屻�?�鍠婇崡鐐差潻闂佸憡锚閻°劑骞堥妸锔剧瘈闁告洦鍘肩粭锟犳⒑閻熸澘妲婚柟铏悾鐑藉Ω閿斿墽鐦堥梺鍛婂姂閸斿本绔熷鍥╃＝闁稿本鑹鹃埀顒勵棑缁牊绗熼�?顒勶�??锟介弽顓炵妞ゆ挾鍣ラ崑銊モ攽椤�?枻渚涢柛鎾寸洴�?�娊鏁冮崒娑氬帾闂婎偄娲㈤崕宕囧閹稿簺浜滈柍鍝勫暙閸樻挳鏌熼绛嬫疁闁轰焦鍔栭幆鏂库攽閸喐娅﹂梻鍌欑劍鐎笛呯矙閹烘鍎庢い鏍ㄥ嚬濞兼牠鏌ц箛姘兼綈鐎规洖顦甸弻鏇熺箾閸喖濮曢梺璇茬箣閻掞妇鎹㈠┑鍡忔灁闁割煈鍠楅悘鎾绘⒑鏉炴壆顦︽い顓犲厴閻涱噣宕�?鑺ユ闂佺粯枪鐏忔瑩藝閵娿儺娓婚柕鍫濇閳锋帡鏌￠崪浣镐喊鐎规洏鍨藉畷锟犳倷閳哄�?�鏉搁梻浣虹帛椤洨鍒掗姘ｆ鐟滃孩绌辨繝鍥舵晝闁挎繂瀛╅悿浣割渻閵堝啫鐏俊顐㈠暣閵嗕線寮崼婵嬪敹闂佺粯鏌ㄩ幖顐︾嵁閸儲鈷掑ù锝囨�?椤曟粎绱掔拠璇ф嫹?閿熶粙鐛繝鍥х疀妞ゆ柨澧介悡瀣攽閻愬弶鈻曞ù婊勭箞閺佹捇鏁撻敓锟??????闂佽鍑界紞鍡涘礈濞戙垺鏅柣鏂垮悑閳锋垿姊洪銈呬粶闁兼椿鍨遍弲鍫曞礈瑜忕壕濂告煕濞嗗浚妲归柕鍥ㄧ箘閳ь剚顔栭崰妤勩亹閸愵喖鐓橀柟杈剧畱闁卞洭鏌曡箛瀣仼缂佺姷鏁诲缁樻媴閸涘﹥鍎撻梺鍝ュ櫏閸嬪﹪骞冭缁绘繈宕堕妸銉ょ暗婵犵數鍋為崹鍫曞春閸愵喖纾婚柟鎹愵嚙�???鍌氼熆鐠虹尨姊楀瑙勬礋濮婄粯绗熸繝鍐�??闂佽法鍠曞Λ鍕嚐椤栨稒娅犻弶鍫㈠亾閿燂拷??闂佽法鍠曟慨銈吤洪幋�???�???闁告劕妯婇崵鏇灻归悩宸剾闁轰礁娲弻锝呂熼崹顔炬闂侀潧鐗炵粻鎾愁潖缂佹ɑ濯村�?�姘煎灡閺侇垶姊虹憴鍕仧濞存粎鍋熼崚鎺撶節濮橆剛顓洪梺缁樏敓�????缂佹顦埞鎴︽倷閺夋垹浠ч梺鎼炲妽濡炰粙宕哄☉銏犵婵°�?�鑳堕崢鍗烆渻閵堝棗濮傞柛濠冩礋瀵悂寮�?崼鐔哄帗濡炪倖鐗楃粙鎺旂矆閸愵喗鐓忛柛銉戝喚浼冮悗娈垮櫘閸撶喎鐣疯ぐ鎺濇晪闁告侗鍓涘Λ顖滅磽閸屾熬�????閿熶粙鎳楅崜浣稿灊妞ゆ牗绮嶅畷鏌ユ煕閺囥劌鐏犵紒鎰殔閳规垿鎮╅煫顓℃姉闂佺粯妫�?鏍惞閸︻厾锛滃┑鈽嗗灥閸嬫劖鏅ラ梻鍌氾拷?锟介崐鎼佸磹閻戣姤鏅搁柨鐕傛�???濠碉紕鍋戦崐鏍垂閻㈢ǹ绠犳慨妞诲亾闁绘侗鍠楃换婵嬪磼閵堝棗缂撻梻渚婃�??閿熻棄鑻晶顔姐亜閺囶亞绉い銏℃礋閺佹捇鏁撻敓�?????缂備讲鍋撻柛鎰ㄦ杺娴滄粓鏌￠崘顭掓嫹?閿熶粙骞忛埄鍐闁绘挸鍑介煬顒佹叏婵犲啯銇濇俊顐㈠暙閳藉顫濋澶嬫瘒闂傚倷鑳堕�?�濠傗枍閺囥垹绠查柛銉墰�?�撲焦淇婇妶鍛櫣闁告濞婇弻鏇＄疀婵犲喛锟???閿熶粙鏌熼柨瀣仢婵﹥妞藉畷銊︾節閸曨厾鏆ら梺璇插閸戝綊宕ｉ崘銊ф殾闁圭儤顨呮儫闂佸啿鎼崐濠氬储闁秵鈷戦梻鍫熻儐瑜版帒纾匡�??锟芥洖娲ㄩ惌鎾寸箾�?�割喕绨奸柣鎾寸洴閹﹢鎮欓悽鍨啒闂佺ǹ瀛╁Λ鎴﹀箯閿燂拷??闂佽法鍠曟慨銈吤洪弽顓熷亯闁稿繘妫跨换鍡樻叏濠靛棛鐒炬俊鏌ョ畺濮婄儤瀵煎▎鎴犳殸闂佺粯顨嗛幐鎼侊綖韫囨梻�???婵﹩鍓涢敍婊冣攽椤旂煫顏勭暦椤掑嫭鏅搁柨鐕傛嫹?缂傚倸鍊搁崐椋庣矆閿燂拷?椤㈡牠宕卞▎鎰闂佺粯鍔欏褔宕瑰┑鍡忔斀闁绘ê寮堕幖鎰版煟閹惧娲撮柡灞剧〒娴狅箓宕滆閸ｎ喚绱撴担鍝勑ｉ柤褰掔畺閳ユ棃宕�?鍢壯囨煕閳╁喚娈旀い顐㈡喘濮婅櫣绮欓崠鈩冩暰濠电偛寮堕…鍥╁垝鐎ｎ喖绠抽柟瀛樻煥閻楁岸姊洪崨濠冪５闁哄懏鐟ч懞杈╂嫚瀹割喗�?�岄梺闈涚墕閹虫劗绮绘导瀛橈�??锟芥慨妯煎帶婢ц揪�????閿熺瓔鍠楁繛濠囧极閹版澘宸濇い蹇撴噺閺夋悂姊绘担鍝勪缓闁稿氦浜竟鏇㈩敇閵忕姵锟??????闂備礁鎼ú锕傛晪婵犳鍠栭崐褰掑Φ閸曨垰顫呴柨娑樺閿燂拷??闂備胶顢婇崑鎰偘閵夆晛�?堟繝闈涱儏濮瑰弶銇勮箛鎾跺闁抽攱甯￠弫鎾绘晸閿燂拷??????闂傚倷鑳堕崢褔宕幐搴㈡珷閹兼番鍔岀粈鍡涙煙閻戞﹩娈㈤柡浣哥Ч閺岋綁骞囬鐔虹▏婵炲瓨绮撴禍璺侯潖濞差亜浼犻柛鏇ㄥ墮閸嬪秹姊洪幖鐐插闁硅櫕鎸哥叅闁秆勵殕閳锋帒霉閿濆懏鎲哥紒澶屽劋娣囧﹪顢曢�?鈥充淮闂佽鍠氶崑銈夊极閸愵喖纾兼慨妯诲敾缁辫鲸绻濆▓鍨灍闁靛洦鐩畷鎴﹀箻缂佹鍘搁柣蹇曞仩椤曆勬叏閸岀偞鐓欐い鏂挎惈閳ь剚绻傞悾鐑藉箳閹存梹�???????闂傚倸鍊峰ù鍥敋瑜忛�?顒佺▓閺呯娀銆佸▎鎾冲唨妞ゆ挾鍋熼悰銉╂⒑閸濆嫭宸濆┑顔芥尦瀹曠懓鈹戦崶鈺冾啎闂佺硶鍓濊摫閻忓浚浜弻宥堫檨闁稿繑绋撳▎銏狀潩椤掑娈ㄩ梺鍦檸閸犳牠锝為崨瀛樼厓闁靛鍎辩敮鐘电磼閵娿儺鐓兼慨濠勭帛閹峰懘宕崟顏勵棜闂備胶鍘х紞濠勭不閺嵮呮殾闁圭増婢樼粻褰掓煥閻曞�?�锟???婵犮垼娉涢オ鏉戭焽閳哄�?�浜滈柟鎹愭硾鍟搁梺浼欑畱閻楁挸顫忛崫鍕懷囧炊瑜忔导鍫濃攽閻愭澘灏冮柛鏇ㄥ弾濞村嫰姊洪幐搴㈢闁稿﹤缍婇幃锟犲即閵忥紕鍘繝鐢靛仜閻忔繈宕濋妶澶嬬厱闁冲搫顑囩粙濠氭煏閸パ冾伃濠殿喒鍋撻梺鏂ユ櫅閸熺�?骞忚ぐ鎺撶厽閹兼番鍔嶅☉褔鏌曢崼鈶跺綊顢氶敐澶婇唶闁哄洨鍋熼敓锟?????闂備礁鎲￠懝楣冨箠韫囨洘宕叉繛鎴炵懄缂嶅洭鏌涢幘�???鍟悡鍌滅磽閸屾瑧顦︽い锕傛涧椤洩顦规い銏″哺婵＄兘鍩℃担渚Ч婵＄偑鍊栭悧�???顫濋妸鈺傛櫢闁跨噦锟???婵犵绱曢崑鎴﹀磹閺嶎偅鏆滈柟铏瑰仦閿燂�???闂佽法鍠撻悺鏃堝礈閻斿鍤曟い鎰╁劘娴滃綊鏌熼悜妯诲皑闁归绮换娑㈠箻閺夋垹鍔伴梺绋款儐閹歌崵鎹㈠☉娆愬�?�闁告劕寮堕惁浠嬫煏婵炵偓娅呴柣鎺炴�???闂備礁鐤囬～澶愬垂閸ф鍨傚Δ锝呭暞閹偞銇勯幇鈺佺仾闁诲繐閰ｉ弻锝嗘償閵堝孩缍堝┑鐐村絻缁绘ê鐣疯ぐ鎺撳癄濠㈣泛鏈▓楣冩⒑闂堟稈搴峰┑鈥虫喘閺佹捇鏁撻敓锟????闂傚倷绀�?幉鈥趁洪敃鍌氱煑閹兼番鍔岄悿�???骞栧ǎ�???濡介柍閿嬪灴閺屾稑鈹戦崱妤婁紝濠碉拷?锟藉级閹�?�寮婚敐澶嬫櫢闁跨噦�????濠碘槅鍋呴悷鈺侇嚕閺屻儱閱囬柡鍥╁枎閿燂�????闂備焦妞块崢浠嬪箰婵犳艾桅闁告洦鍨扮粻绛规嫹?閿熷鍎遍ˇ浼搭敁閺嶃劎绠鹃悗娑欘焽閻绱掗鑲┬у┑锛勬暬�?�曠喖顢涘杈╂澑闂備礁鐤囧銊╂嚄閸洖绀夐柡澶嬪灍锟??浠嬫煃閵夈儱鏆辩紒鐙欏洦鐓欐い鏃傚帶閳ь剙鐏濋锝嗙節濮橆厽娅滄繝銏ｆ硾椤戝棗鈻嶅⿰鍫熲拺闁告稑锕ｇ欢閬嶆煕濡鐏婄紒銊︽そ濮婂宕掑▎鎰垫▊缂備線纭搁崰姘嚗婵犲洤绀堢憸搴＄暦閺屻儲鐓曟い鎰剁悼缁犳﹢鏌￠崱顓犵暤闁哄矉缍佸锟??宕掑Δ浣哥彵闂備浇妗ㄧ粈浣肝涘┑�?�摕婵炴垶鐭▽顏堟煙鐟欏嫬濮囨い銉︾箘缁辨挻鎷呴崫鍕戠偤鏌涙惔銊︽锭妞ゎ偄绻戠换婵嗩潩椤掑偊绱叉繝鐢靛仜濡瑩宕归崹顐＄箚濞寸姴顑嗛埛鎴犵磼鐎ｎ亝鍋ユい搴㈩殜閺屾盯鎮㈤柨�?�淮濠电姭鍋撳ù锝囩《锟??鑺ャ亜閺冨浂娼￠柣鐔稿閺嬫牗绻涢幋鐐跺妞ゃ儲姘ㄩ幉鎼佹偋閸繄鐟查梺绋匡功閺佸寮婚妸銉㈡斀闁糕剝渚楅埀顒侇殕缁绘盯宕ㄩ鍡嫹?閿熶粙鏌＄仦绋垮⒉闁瑰嚖�???????闂傚倷绀�?幖顐�?嫉椤掑嫭鍎庢い鏍亼閳ь兛绶氬鎾閳哄倹娅囬梻�???娼х换鎺撳垔椤撶儐鐒介柛鎾�?懐锛濋梺绋挎湰閻熝囁囬敂濮愪簻闁瑰瓨绻冮崳浠嬫煙楠炲灝鐏叉鐐叉喘�?�墎鎹勯妸銉ョ闂傚�?�鑳堕�?�濠囧箵椤忓牊鈷旈柛鏇ㄥ灠绾惧鏌熼柇锟??鏋ょ痪鎹愭闇夐柨婵嗙墕娴滄鏌熸潏楣冩闁绘挶鍎查妵鍕箻鐠哄搫澹夊┑鐐存尭椤兘寮婚弴銏犻唶婵犻潧娴傚Λ鐐烘⒑鐠囪尙绠為柛搴ｆ暬�?�鎮㈤崗鍏煎劒濡炪�?�鍔戦崹褰掞綖锟??鍕拺閻庡湱濮甸ˉ澶嬨亜閿旂偓鏆鐐插暣閹儳鐣濋埀顒勬儗濞嗘挻鍋ｉ柟顓熷笒婵＄厧鈹戦鍡涙濞ｅ洤锕幃娆擃敂鎼淬垹锟???闂佽法鍠撻弲顐﹀极閿燂拷?閺佹捇鏁撻敓�??????濠殿喗顭囬崢褍顕ｉ敓�????閺屾盯鍩￠崒婊勫垱濡ょ姷鍋涢澶愬箖閳哄懏鍋ㄧ痪鏉款槺闂傤垱绻濋悽闈涗哗闁规椿浜炲濠冪鐎ｅ墎绋忛梺鍝勭▉閸欏酣寮崒鐐寸厱婵炴垵宕弸娑虫嫹?閿熺瓔鍠栧鈥愁潖濞差亜绠归柣鎰絻婵爼姊洪崨濠冨鞍閿燂拷?閹间礁绠栭柨鐔哄У閸嬪嫰鏌ゅù�?�珔鐟滄澘瀚板娲箹閻愭彃濮岄梺鍛婃煥缁夊綊骞冮敓鐘参ㄩ柍鍝勶拷?锟介崢鍗炩攽閻樼粯娑ч柣锟??妫濆畷婵撴嫹?閿熺瓔鍠楅悡蹇涙煕閵夋垵鍠氶敓锟?????闂傚倷鐒﹂崜姘跺储閹间礁鐤炬繝濠傜墕閸ㄥ倻鎲搁悧鍫濈瑨缂佺姵鐓￠弻鏇＄疀閺囩倫娑㈡煛閳ь剚绂掞�??锟筋偆鍘遍梺璺ㄥ櫐閿燂拷??闂佸搫鎳忕划鎾崇暦閹剧粯顥堟繛鎴ｉ哺鐎靛矂姊洪棃娑氬婵☆偅鐟ф禍鎼佸箥椤斿墽锛滈柣搴秵閸嬪嫮绮閺屽秷顧�?柛鎾寸缁岄亶宕崟搴㈢洴�?�曠喖顢涘鍗炲箣闂備胶顢婇幓顏堟⒔閸曨垰纾归柣鎴ｅГ閻撶�?鏌熼梻�?�稿妽婵炴嚪鍕闁瑰啿鍢查幊鎰閽樺褰掓晲閸ャ劌娈�?紓浣藉皺缁垳鎹㈤敓�????????闂備椒绱徊鍧楀礂濡警鍤曢柟缁㈠枛椤懘鏌ｅΟ鑽ゅ灩闁告劕澧介崬鐢告煟閻樼儤顏犻悘蹇嬪妼椤斿繘濡烽埡鍌滃幍濡炪�?�鐗楃划灞剧鏉堛劍鍙忓┑鐘插暞閵囨繈鏌＄仦鑺ュ殗闁诡喗鐟╅幊鐘垫崉娓氼垯绱�?繝鐢靛Л閹峰啴宕橀鍛枛闂備緤锟???閿熺晫鈹掗柛鏂跨Ф閹广垹鈹戯拷?锟筋亞顦ㄩ梺宕囨�?閵囨﹢鎼规惔顫箚闁靛牆娲ゅ暩闂佺ǹ顑囬崑銈夊箖瑜旈幃鈺冩嫚閼碱剛鏆繝鐢靛Т閿曘�?�鎮ч崱娑欙拷?锟藉┑鐘叉处閻撳繐鈹戦悙鑼虎闁告梹鎸抽弫鎾绘晸閿燂�?????闂傚倸鍊搁崐鎼佸磹�?�勬噴褰掑炊瑜夐弸鏍煛閸ャ儱鐏╃紒鎰殘閳ь剙绠嶉崕鍗灻洪妶澶婂瀭婵犻潧娲ㄧ粻楣冩煕閳╁叐鎴犱焊椤撶姷纾奸柣妯虹－婢ч亶鏌熼崣澶嬶�??锟斤�??锟筋噮鍣ｅ畷鐓庘攽閸垺姣囬梻鍌欑閸熷潡骞栭�???鐤い鏍ワ拷?锟介敓锟????闂佽法鍠曟慨銈呯暆閹间礁钃熸繛鎴炃氶弸搴ㄧ叓閸ラ绋诲Δ鏃堟⒒閿燂�??閳ь剛鍋涢懟顖涙櫠婵犳碍鐓曢柟鎹愭硾閺嬪孩銇勯銏㈢閻撱倖銇勮箛鎾村櫣濞寸媭鍙冨娲传閸曞灚笑缂備降鍔戞禍鍫曠嵁閹版澘�?冩い蹇撴閿涙繃绻涢幘纾嬪婵炲眰鍊曢埢宥咁潨閳ь剟寮诲☉銏犖╅柕濠忓閵嗘劕顪冮妶鍡樼┛缂傚秳绀�?锝嗙節濮橆儵銊╂煏婢诡垰鑻弲锝嗙�?閻㈤潧浠╅柟娲讳簽�?�板﹪鎸婃径娑虫�??閿熶粙姊洪敓�????缁夋挳鎯屽Δ鍛厱闁斥晛鍟伴埊鏇㈡煃闁垮鐏╃紒杈ㄦ尰閹峰懘鎯傞崨濠傤�????闂傚倸鍊烽懗鑸电仚闂佹寧娲忛崐鏇㈡晝閵忋倖鐒硷拷?锟姐儱鎳愰崝�???顪冮妶鍡楃瑐闁煎啿鐖煎畷顖炲蓟閵夛妇�??????
        .axi_wen_o(axi_wen),
        .axi_waddr_o(axi_waddr),
        .axi_wdata_o(axi_wdata),
        .axi_wvalid_o(axi_wvalid),
        .axi_wlast_o(axi_wlast),
        .axi_wlen_o(axi_wlen)
    );


`ifdef DIFF
        wire [31:0] debug_wb_pc_diff0       ;
        wire [31:0] debug_wb_inst_diff0     ;
        wire [3:0]  debug_wb_rf_wen_diff0   ;
        wire [4:0]  debug_wb_rf_wnum_diff0  ;
        wire [31:0] debug_wb_rf_wdata_diff0 ;

        wire [31:0] debug_wb_pc_diff1       ;
        wire [31:0] debug_wb_inst_diff1     ;
        wire [ 3:0] debug_wb_rf_wen_diff1   ;
        wire [ 4:0] debug_wb_rf_wnum_diff1  ;
        wire [31:0] debug_wb_rf_wdata_diff1 ;

        wire        inst_valid_diff0        ;
        wire        cnt_inst_diff0          ;
        wire        csr_rstat_en_diff0      ;
        wire [31:0] csr_data_diff0          ;

        wire        inst_valid_diff1        ;
        wire        cnt_inst_diff1          ;
        wire        csr_rstat_en_diff1      ;
        wire [31:0] csr_data_diff1          ;

        wire        excp_flush_diff0        ;
        wire        ertn_flush_diff0        ;
        wire [ 5:0] ecode_diff0             ;

        wire        excp_flush_diff1        ;
        wire        ertn_flush_diff1        ;
        wire [ 5:0] ecode_diff1             ;

        wire [ 7:0] inst_st_en_diff0        ;
        wire [31:0] st_paddr_diff0          ;
        wire [31:0] st_vaddr_diff0          ;
        wire [31:0] st_data_diff0           ;

        wire [ 7:0] inst_st_en_diff1        ;
        wire [31:0] st_paddr_diff1          ;
        wire [31:0] st_vaddr_diff1          ;
        wire [31:0] st_data_diff1           ;

        wire [ 7:0] inst_ld_en_diff0        ;
        wire [31:0] ld_paddr_diff0          ;
        wire [31:0] ld_vaddr_diff0          ;

        wire [ 7:0] inst_ld_en_diff1        ;
        wire [31:0] ld_paddr_diff1          ;
        wire [31:0] ld_vaddr_diff1          ;

        wire        tlbfill_en_diff0        ;
        wire        tlbfill_en_diff1        ;

        assign {    debug_wb_pc_diff0,
                    debug_wb_inst_diff0,
                    debug_wb_rf_wen_diff0,
                    debug_wb_rf_wnum_diff0,
                    debug_wb_rf_wdata_diff0,

                    inst_valid_diff0,
                    cnt_inst_diff0,
                    csr_rstat_en_diff0,
                    csr_data_diff0,

                    excp_flush_diff0,
                    ertn_flush_diff0,
                    ecode_diff0,

                    inst_st_en_diff0,
                    st_paddr_diff0,
                    st_vaddr_diff0,
                    st_data_diff0,

                    inst_ld_en_diff0,
                    ld_paddr_diff0,
                    ld_vaddr_diff0,

                    tlbfill_en_diff0} = diff0;

        assign {    debug_wb_pc_diff1,
                    debug_wb_inst_diff1,
                    debug_wb_rf_wen_diff1,
                    debug_wb_rf_wnum_diff1,
                    debug_wb_rf_wdata_diff1,

                    inst_valid_diff1,
                    cnt_inst_diff1,
                    csr_rstat_en_diff1,
                    csr_data_diff1,

                    excp_flush_diff1,
                    ertn_flush_diff1,
                    ecode_diff1,

                    inst_st_en_diff1,
                    st_paddr_diff1,
                    st_vaddr_diff1,
                    st_data_diff1,

                    inst_ld_en_diff1,
                    ld_paddr_diff1,
                    ld_vaddr_diff1,

                    tlbfill_en_diff1} = diff1;

    always @(posedge aclk) begin
        if (rst) begin
            {cmt0_valid, cmt0_cnt_inst, cmt0_timer_64, cmt0_inst_ld_en, cmt0_ld_paddr, cmt0_ld_vaddr, cmt0_inst_st_en, cmt0_st_paddr, cmt0_st_vaddr, cmt0_st_data, cmt0_csr_rstat_en, cmt0_csr_data} <= 0;
            {cmt0_wen, cmt0_wdest, cmt0_wdata, cmt0_pc, cmt0_inst} <= 0;
            {trap, trap_code, cycleCnt, instrCnt} <= 0;
        end
        else begin
            cmt0_valid       <= inst_valid_diff0;
            cmt0_cnt_inst    <= cnt_inst_diff0;
            cmt0_timer_64    <= cnt;
            cmt0_inst_ld_en  <= inst_ld_en_diff0;
            cmt0_ld_paddr    <= ld_paddr_diff0;
            cmt0_ld_vaddr    <= ld_vaddr_diff0;
            cmt0_inst_st_en  <= inst_st_en_diff0;
            cmt0_st_paddr    <= st_paddr_diff0;
            cmt0_st_vaddr    <= st_vaddr_diff0;
            cmt0_st_data     <= st_data_diff0;
            cmt0_csr_rstat_en<= csr_rstat_en_diff0;
            cmt0_csr_data    <= csr_data_diff0;

            cmt0_wen         <= debug_wb_rf_wen_diff0;
            cmt0_wdest       <= {3'd0, debug_wb_rf_wnum_diff0};

            cmt0_wdata       <= debug_wb_rf_wdata_diff0;
            cmt0_pc          <= debug_wb_pc_diff0;
            cmt0_inst        <= debug_wb_inst_diff0;

            cmt0_excp_flush  <= excp_flush_diff0;
            cmt0_ertn        <= ertn_flush_diff0;
            cmt0_csr_ecode   <= ecode_diff0;
            cmt0_tlbfill_en  <= tlbfill_en_diff0;   

            cmt1_valid       <= inst_valid_diff1;
            cmt1_cnt_inst    <= cnt_inst_diff1;
            cmt1_timer_64    <= cnt;
            cmt1_inst_ld_en  <= inst_ld_en_diff1;
            cmt1_ld_paddr    <= ld_paddr_diff1;
            cmt1_ld_vaddr    <= ld_vaddr_diff1;
            cmt1_inst_st_en  <= inst_st_en_diff1;
            cmt1_st_paddr    <= st_paddr_diff1;
            cmt1_st_vaddr    <= st_vaddr_diff1;
            cmt1_st_data     <= st_data_diff1;
            cmt1_csr_rstat_en<= csr_rstat_en_diff1;
            cmt1_csr_data    <= csr_data_diff1;

            cmt1_wen         <= debug_wb_rf_wen_diff1;
            cmt1_wdest       <= {3'd0, debug_wb_rf_wnum_diff1};

            cmt1_wdata       <= debug_wb_rf_wdata_diff1;
            cmt1_pc          <= debug_wb_pc_diff1;
            cmt1_inst        <= debug_wb_inst_diff1;

            cmt1_excp_flush  <= excp_flush_diff1;
            cmt1_ertn        <= ertn_flush_diff1;
            cmt1_csr_ecode   <= ecode_diff1;
            cmt1_tlbfill_en  <= tlbfill_en_diff1;
            cmt_rand_index   <= cnt[4:0];  

            regs_diff        <= regs_diff_out;
        end
          
    end

    assign debug0_wb_inst = debug_wb_inst_diff0;
    assign debug0_wb_pc = debug_wb_pc_diff0;
    assign debug0_wb_rf_wen = debug_wb_rf_wen_diff0;
    assign debug0_wb_rf_wnum = debug_wb_rf_wnum_diff0;
    assign debug0_wb_rf_wdata = debug_wb_rf_wdata_diff0;

    assign debug1_wb_inst = debug_wb_inst_diff1;
    assign debug1_wb_pc = debug_wb_pc_diff1;
    assign debug1_wb_rf_wen = debug_wb_rf_wen_diff1;
    assign debug1_wb_rf_wnum = debug_wb_rf_wnum_diff1;
    assign debug1_wb_rf_wdata = debug_wb_rf_wdata_diff1;

    assign debug_wb_pc       = debug0_wb_pc      | debug1_wb_pc      ;
    assign debug_wb_rf_we    = debug0_wb_rf_wen  | debug1_wb_rf_wen  ;
    assign debug_wb_rf_wnum  = debug0_wb_rf_wnum | debug1_wb_rf_wnum ;
    assign debug_wb_rf_wdata = debug0_wb_rf_wdata| debug1_wb_rf_wdata;



    reg [63:0] inst_num;
    always @( posedge aclk ) begin
        if (rst) begin
            inst_num <= 0;
        end else if (inst_valid_diff0 && inst_valid_diff1) begin
            inst_num <= inst_num + 2;
        end else if (inst_valid_diff0 || inst_valid_diff1) begin
            inst_num <= inst_num + 1;
        end else begin
            inst_num <= inst_num;
        end
    end

    always @(posedge aclk) begin
        if (rst) begin
            {trap, trap_code, cycleCnt, instrCnt} <= 0;
        end else begin
            trap            <= 0                        ;
            trap_code       <= regs_diff[10][7:0]       ;
            cycleCnt        <= cycleCnt + 1             ;
            instrCnt        <= instrCnt;
        end
    end

    reg excp_flush;
    reg [31:0] excp_pc;
    reg [31:0] excp_inst;
    
    always @(*) begin
        if (cmt0_excp_flush) begin
            excp_flush = cmt0_excp_flush;
            excp_pc = cmt0_pc;
            excp_inst = cmt0_inst;
        end else begin
            excp_flush = cmt1_excp_flush;
            excp_pc = cmt1_pc;
            excp_inst = cmt1_inst;
        end
    end

    DifftestInstrCommit DifftestInstrCommit_0(
        .clock              (aclk           ),
        .coreid             (0              ),
        .index              (0     ),
        .valid              (cmt0_valid   ),
        .pc                 (cmt0_pc      ),
        .instr              (cmt0_inst    ),
        .skip               (0              ),
        .is_TLBFILL         (cmt0_tlbfill_en),
        .TLBFILL_index      (cmt_rand_index ),
        .is_CNTinst         (cmt0_cnt_inst),
        .timer_64_value     (cmt0_timer_64),
        .wen                (cmt0_wen     ),
        .wdest              (cmt0_wdest   ),
        .wdata              (cmt0_wdata   ),
        .csr_rstat          (cmt0_csr_rstat_en),
        .csr_data           (cmt0_csr_data)
    );

    DifftestInstrCommit DifftestInstrCommit_1(
        .clock              (aclk           ),
        .coreid             (0              ),
        .index              (1    ),
        .valid              (cmt1_valid   ),
        .pc                 (cmt1_pc      ),
        .instr              (cmt1_inst    ),
        .skip               (0              ),
        .is_TLBFILL         (cmt1_tlbfill_en),
        .TLBFILL_index      (cmt_rand_index ),
        .is_CNTinst         (cmt1_cnt_inst),
        .timer_64_value     (cmt1_timer_64),
        .wen                (cmt1_wen     ),
        .wdest              (cmt1_wdest   ),
        .wdata              (cmt1_wdata   ),
        .csr_rstat          (cmt1_csr_rstat_en),
        .csr_data           (cmt1_csr_data)
    );



    DifftestExcpEvent DifftestExcpEvent(
        .clock              (aclk           ),
        .coreid             (0              ),
        .excp_valid         (excp_flush     ),
        .eret               (cmt0_ertn      ),
        .intrNo             (csr_estat_diff_0[12:2]),
        .cause              (cmt0_csr_ecode ),
        .exceptionPC        (excp_pc        ),
        .exceptionInst      (excp_inst      )
    );

    DifftestTrapEvent DifftestTrapEvent(
        .clock              (aclk           ),
        .coreid             (0              ),
        .valid              (trap           ),
        .code               (trap_code      ),
        .pc                 (cmt0_pc        ),
        .cycleCnt           (cycleCnt       ),
        .instrCnt           (instrCnt       )
    );
     
    DifftestStoreEvent DifftestStoreEvent0(
        .clock              (aclk             ),
        .coreid             (0                ),
        .index              (0                ),
        .valid              (cmt0_inst_st_en),
        .storePAddr         (cmt0_st_paddr  ),
        .storeVAddr         (cmt0_st_vaddr  ),
        .storeData          (cmt0_st_data   )
    );

    DifftestStoreEvent DifftestStoreEvent1(
        .clock              (aclk             ),
        .coreid             (0                ),
        .index              (1                ),
        .valid              (cmt1_inst_st_en),
        .storePAddr         (cmt1_st_paddr  ),
        .storeVAddr         (cmt1_st_vaddr  ),
        .storeData          (cmt1_st_data   )
    );

    DifftestLoadEvent DifftestLoadEvent0(
        .clock              (aclk             ),
        .coreid             (0                ),
        .index              (0                ),
        .valid              (cmt0_inst_ld_en),
        .paddr              (cmt0_ld_paddr  ),
        .vaddr              (cmt0_ld_vaddr  )
    );

    DifftestLoadEvent DifftestLoadEvent1(
        .clock              (aclk             ),
        .coreid             (0                ),
        .index              (1                ),
        .valid              (cmt1_inst_ld_en),
        .paddr              (cmt1_ld_paddr  ),
        .vaddr              (cmt1_ld_vaddr  )
    );

    DifftestCSRRegState DifftestCSRRegState(
        .clock              (aclk               ),
        .coreid             (0                  ),
        .crmd               (csr_crmd_diff_0    ),
        .prmd               (csr_prmd_diff_0    ),
        .euen               (0                  ),
        .ecfg               (csr_ectl_diff_0    ),
        .estat              (csr_estat_diff_0   ),
        .era                (csr_era_diff_0     ),
        .badv               (csr_badv_diff_0    ),
        .eentry             (csr_eentry_diff_0  ),
        .tlbidx             (csr_tlbidx_diff_0  ),
        .tlbehi             (csr_tlbehi_diff_0  ),
        .tlbelo0            (csr_tlbelo0_diff_0 ),
        .tlbelo1            (csr_tlbelo1_diff_0 ),
        .asid               (csr_asid_diff_0    ),
        .pgdl               (csr_pgdl_diff_0    ),
        .pgdh               (csr_pgdh_diff_0    ),
        .save0              (csr_save0_diff_0   ),
        .save1              (csr_save1_diff_0   ),
        .save2              (csr_save2_diff_0   ),
        .save3              (csr_save3_diff_0   ),
        .tid                (csr_tid_diff_0     ),
        .tcfg               (csr_tcfg_diff_0    ),
        .tval               (csr_tval_diff_0    ),
        .ticlr              (csr_ticlr_diff_0   ),
        .llbctl             (csr_llbctl_diff_0  ),
        .tlbrentry          (csr_tlbrentry_diff_0),
        .dmw0               (csr_dmw0_diff_0    ),
        .dmw1               (csr_dmw1_diff_0    )
    );

    DifftestGRegState DifftestGRegState(
        .clock              (aclk       ),
        .coreid             (0          ),
        .gpr_0              (0          ),
        .gpr_1              (regs_diff[1]   ),
        .gpr_2              (regs_diff[2]   ),
        .gpr_3              (regs_diff[3]   ),
        .gpr_4              (regs_diff[4]   ),
        .gpr_5              (regs_diff[5]   ),
        .gpr_6              (regs_diff[6]   ),
        .gpr_7              (regs_diff[7]   ),
        .gpr_8              (regs_diff[8]   ),
        .gpr_9              (regs_diff[9]   ),
        .gpr_10             (regs_diff[10]   ),
        .gpr_11             (regs_diff[11]   ),
        .gpr_12             (regs_diff[12]   ),
        .gpr_13             (regs_diff[13]   ),
        .gpr_14             (regs_diff[14]   ),
        .gpr_15             (regs_diff[15]   ),
        .gpr_16             (regs_diff[16]   ),
        .gpr_17             (regs_diff[17]   ),
        .gpr_18             (regs_diff[18]   ),
        .gpr_19             (regs_diff[19]   ),
        .gpr_20             (regs_diff[20]   ),
        .gpr_21             (regs_diff[21]   ),
        .gpr_22             (regs_diff[22]   ),
        .gpr_23             (regs_diff[23]   ),
        .gpr_24             (regs_diff[24]   ),
        .gpr_25             (regs_diff[25]   ),
        .gpr_26             (regs_diff[26]   ),
        .gpr_27             (regs_diff[27]   ),
        .gpr_28             (regs_diff[28]   ),
        .gpr_29             (regs_diff[29]   ),
        .gpr_30             (regs_diff[30]   ),
        .gpr_31             (regs_diff[31]   )
    );
    
    
    `endif

/*
    wire [101:0] data1;
    wire [101:0] data2;
    wire valid1;
    wire valid2;
    wire [101:0] debug_data_out;
    wire debug_valid_out;

    assign data1 = {debug_wb_we1,debug_reg_addr1,debug_wdata1,debug_inst1,debug_pc1};
    assign data2 = {debug_wb_we2,debug_reg_addr2,debug_wdata2,debug_inst2,debug_pc2};
    assign valid1 = debug_wb_valid1;
    assign valid2 = debug_wb_valid2;

    debug_FIFO debug
    (
        .clk(aclk),
        .rst(rst),
        .valid1(valid1),
        .data1(data1),
        .valid2(valid2),
        .data2(data2),
        .data_out(debug_data_out),
        .valid_out(debug_valid_out)
    );

    assign debug0_wb_pc = debug_data_out[31:0];  
    assign debug0_wb_rf_wen = {4{debug_data_out[101]}};
    assign debug0_wb_rf_wnum = debug_data_out[100:96];
    assign debug0_wb_rf_wdata = debug_data_out[95:64];
*/



endmodule