`ifndef CSR_DEFINES_V
`define CSR_DEFINES_V

// CSR 地址
`define CSR_CRMD        14'b00000000000000  //0
`define CSR_PRMD        14'b00000000000001  //1
`define CSR_EUEN        14'b00000000000010  //2
`define CSR_ECFG        14'b00000000000100  //4
`define CSR_ESTAT       14'b00000000000101  //5
`define CSR_ERA         14'b00000000000110  //6
`define CSR_BADV        14'b00000000000111  //7
`define CSR_EENTRY      14'b00000000001100  //c
`define CSR_TLBIDX      14'b00000000010000  //10
`define CSR_TLBEHI      14'b00000000010001  //11
`define CSR_TLBELO0     14'b00000000010010  //12
`define CSR_TLBELO1     14'b00000000010011  //13
`define CSR_ASID        14'b00000000011000  //18
`define CSR_PGDL        14'b00000000011001  //19
`define CSR_PGDH        14'b00000000011010  //1a
`define CSR_PGD         14'b00000000011011  //1b
`define CSR_CPUID       14'b00000000100000  //20
`define CSR_SAVE0       14'b00000000110000  //30
`define CSR_SAVE1       14'b00000000110001  //31
`define CSR_SAVE2       14'b00000000110010  //32
`define CSR_SAVE3       14'b00000000110011  //33
`define CSR_TID         14'b00000001000000  //40
`define CSR_TCFG        14'b00000001000001  //41
`define CSR_TVAL        14'b00000001000010  //42
`define CSR_TICLR       14'b00000001000100  //44
`define CSR_LLBCTL      14'b00000001100000  //60
`define CSR_TLBRENTRY   14'b00000010001000  //80
`define CSR_CTAG        14'b00000010011000  //98
`define CSR_DMW0        14'b00000110000000  //180
`define CSR_DMW1        14'b00000110000001  //181
`define CSR_CPUCFG1     14'b00000010110001  
`define CSR_CPUCFG2     14'b00000010110010
`define CSR_CPUCFG10    14'b00000011000000
`define CSR_CPUCFG11    14'b00000011000001
`define CSR_CPUCFG12    14'b00000011000010
`define CSR_CPUCFG13    14'b00000011000011

// Exceptions
`define EXCEPTION_INT 7'b0000000   //0
`define EXCEPTION_PIL 7'b0000010   //2
`define EXCEPTION_PIS 7'b0000100   //4
`define EXCEPTION_PIF 7'b0000110   //6
`define EXCEPTION_PME 7'b0001000   //8
`define EXCEPTION_PPI 7'b0001110   //e
`define EXCEPTION_ADEF 7'b0010000   //10
`define EXCEPTION_ADEM 7'b0010001   //11
`define EXCEPTION_ALE 7'b0010010   //12
`define EXCEPTION_SYS 7'b0010110   //16
`define EXCEPTION_BRK 7'b0011000   //18
`define EXCEPTION_INE 7'b0011010   //1a
`define EXCEPTION_IPE 7'b0011100   //1c
`define EXCEPTION_FPD 7'b0011110   //1e
`define EXCEPTION_FPE 7'b0100100   //24
`define EXCEPTION_TLBR 7'b1111110   //7e
`define EXCEPTION_NOP 7'b1111111   //7f

`endif
